library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------
-- synthesis translate_off 
library ims;
use ims.coprocessor.all;
use ims.conversion.all;
-- synthesis translate_on 
-------------------------------------------------------------------------

ENTITY Q16_8_C_to_V_RAM is
	PORT (
		RESET    : in  STD_LOGIC;
		CLOCK    : in  STD_LOGIC;
		HOLDN    : in  std_ulogic;
		WRITE_EN : in  STD_LOGIC;
		READ_EN  : in  STD_LOGIC;
		INPUT_1  : in  STD_LOGIC_VECTOR(31 downto 0);
		OUTPUT_1 : out STD_LOGIC_VECTOR(31 downto 0)
	);
END;

architecture cRAM of Q16_8_C_to_V_RAM is
   type ram_type is array (0 to 1824-1) of STD_LOGIC_VECTOR (15 downto 0);                 
   type rom_type is array (0 to 1824-1) of UNSIGNED (10 downto 0);                 
   signal RAM : ram_type;

   constant ROM : rom_type:= (
		TO_UNSIGNED(  75, 11), TO_UNSIGNED( 618, 11), TO_UNSIGNED( 732, 11), TO_UNSIGNED(1425, 11), TO_UNSIGNED(1500, 11), TO_UNSIGNED(1683, 11), TO_UNSIGNED(  84, 11), TO_UNSIGNED( 621, 11), 
		TO_UNSIGNED( 738, 11), TO_UNSIGNED(1428, 11), TO_UNSIGNED(1506, 11), TO_UNSIGNED(1614, 11), TO_UNSIGNED(  86, 11), TO_UNSIGNED( 624, 11), TO_UNSIGNED( 744, 11), TO_UNSIGNED(1437, 11), 
		TO_UNSIGNED(1488, 11), TO_UNSIGNED(1819, 11), TO_UNSIGNED(  12, 11), TO_UNSIGNED(  88, 11), TO_UNSIGNED( 627, 11), TO_UNSIGNED( 750, 11), TO_UNSIGNED(1440, 11), TO_UNSIGNED(1512, 11), 
		TO_UNSIGNED(  15, 11), TO_UNSIGNED(  90, 11), TO_UNSIGNED( 630, 11), TO_UNSIGNED( 756, 11), TO_UNSIGNED(1443, 11), TO_UNSIGNED(1524, 11), TO_UNSIGNED(  18, 11), TO_UNSIGNED(  92, 11), 
		TO_UNSIGNED( 633, 11), TO_UNSIGNED( 762, 11), TO_UNSIGNED(1446, 11), TO_UNSIGNED(1518, 11), TO_UNSIGNED(  21, 11), TO_UNSIGNED(  94, 11), TO_UNSIGNED( 636, 11), TO_UNSIGNED( 768, 11), 
		TO_UNSIGNED(1449, 11), TO_UNSIGNED(1542, 11), TO_UNSIGNED(  24, 11), TO_UNSIGNED(  96, 11), TO_UNSIGNED( 639, 11), TO_UNSIGNED( 774, 11), TO_UNSIGNED(1452, 11), TO_UNSIGNED(1548, 11), 
		TO_UNSIGNED(  27, 11), TO_UNSIGNED(  98, 11), TO_UNSIGNED( 642, 11), TO_UNSIGNED( 780, 11), TO_UNSIGNED(1455, 11), TO_UNSIGNED(1530, 11), TO_UNSIGNED(  30, 11), TO_UNSIGNED( 100, 11), 
		TO_UNSIGNED( 645, 11), TO_UNSIGNED( 786, 11), TO_UNSIGNED(1461, 11), TO_UNSIGNED(1536, 11), TO_UNSIGNED(  33, 11), TO_UNSIGNED( 102, 11), TO_UNSIGNED( 648, 11), TO_UNSIGNED( 792, 11), 
		TO_UNSIGNED(1458, 11), TO_UNSIGNED(1554, 11), TO_UNSIGNED(  36, 11), TO_UNSIGNED( 104, 11), TO_UNSIGNED( 651, 11), TO_UNSIGNED( 798, 11), TO_UNSIGNED(1485, 11), TO_UNSIGNED(1560, 11), 
		TO_UNSIGNED(  39, 11), TO_UNSIGNED( 106, 11), TO_UNSIGNED( 654, 11), TO_UNSIGNED( 804, 11), TO_UNSIGNED(1572, 11), TO_UNSIGNED(1617, 11), TO_UNSIGNED(  42, 11), TO_UNSIGNED( 108, 11), 
		TO_UNSIGNED( 657, 11), TO_UNSIGNED( 810, 11), TO_UNSIGNED(1398, 11), TO_UNSIGNED(1566, 11), TO_UNSIGNED(  45, 11), TO_UNSIGNED( 110, 11), TO_UNSIGNED( 660, 11), TO_UNSIGNED( 816, 11), 
		TO_UNSIGNED(1401, 11), TO_UNSIGNED(1584, 11), TO_UNSIGNED(  48, 11), TO_UNSIGNED( 112, 11), TO_UNSIGNED( 663, 11), TO_UNSIGNED( 822, 11), TO_UNSIGNED(1404, 11), TO_UNSIGNED(1578, 11), 
		TO_UNSIGNED(  51, 11), TO_UNSIGNED( 114, 11), TO_UNSIGNED( 666, 11), TO_UNSIGNED( 828, 11), TO_UNSIGNED(1413, 11), TO_UNSIGNED(1596, 11), TO_UNSIGNED(  54, 11), TO_UNSIGNED( 116, 11), 
		TO_UNSIGNED( 669, 11), TO_UNSIGNED( 690, 11), TO_UNSIGNED(1416, 11), TO_UNSIGNED(1602, 11), TO_UNSIGNED(  57, 11), TO_UNSIGNED( 118, 11), TO_UNSIGNED( 672, 11), TO_UNSIGNED( 696, 11), 
		TO_UNSIGNED(1419, 11), TO_UNSIGNED(1590, 11), TO_UNSIGNED(   0, 11), TO_UNSIGNED(  60, 11), TO_UNSIGNED( 120, 11), TO_UNSIGNED( 675, 11), TO_UNSIGNED( 702, 11), TO_UNSIGNED(1407, 11), 
		TO_UNSIGNED(  63, 11), TO_UNSIGNED( 122, 11), TO_UNSIGNED( 678, 11), TO_UNSIGNED( 708, 11), TO_UNSIGNED(1410, 11), TO_UNSIGNED(1476, 11), TO_UNSIGNED(  66, 11), TO_UNSIGNED( 124, 11), 
		TO_UNSIGNED( 681, 11), TO_UNSIGNED( 714, 11), TO_UNSIGNED(1434, 11), TO_UNSIGNED(1464, 11), TO_UNSIGNED(  69, 11), TO_UNSIGNED( 126, 11), TO_UNSIGNED( 684, 11), TO_UNSIGNED( 720, 11), 
		TO_UNSIGNED(1431, 11), TO_UNSIGNED(1470, 11), TO_UNSIGNED(  72, 11), TO_UNSIGNED( 128, 11), TO_UNSIGNED( 687, 11), TO_UNSIGNED( 726, 11), TO_UNSIGNED(1422, 11), TO_UNSIGNED(1494, 11), 
		TO_UNSIGNED( 186, 11), TO_UNSIGNED( 234, 11), TO_UNSIGNED( 775, 11), TO_UNSIGNED( 906, 11), TO_UNSIGNED(1435, 11), TO_UNSIGNED(1585, 11), TO_UNSIGNED( 188, 11), TO_UNSIGNED( 236, 11), 
		TO_UNSIGNED( 781, 11), TO_UNSIGNED( 909, 11), TO_UNSIGNED(1432, 11), TO_UNSIGNED(1579, 11), TO_UNSIGNED( 190, 11), TO_UNSIGNED( 238, 11), TO_UNSIGNED( 787, 11), TO_UNSIGNED( 912, 11), 
		TO_UNSIGNED(1423, 11), TO_UNSIGNED(1597, 11), TO_UNSIGNED( 192, 11), TO_UNSIGNED( 240, 11), TO_UNSIGNED( 793, 11), TO_UNSIGNED( 915, 11), TO_UNSIGNED(1426, 11), TO_UNSIGNED(1603, 11), 
		TO_UNSIGNED( 194, 11), TO_UNSIGNED( 242, 11), TO_UNSIGNED( 799, 11), TO_UNSIGNED( 918, 11), TO_UNSIGNED(1429, 11), TO_UNSIGNED(1591, 11), TO_UNSIGNED(   1, 11), TO_UNSIGNED( 196, 11), 
		TO_UNSIGNED( 244, 11), TO_UNSIGNED( 805, 11), TO_UNSIGNED( 921, 11), TO_UNSIGNED(1438, 11), TO_UNSIGNED( 198, 11), TO_UNSIGNED( 246, 11), TO_UNSIGNED( 811, 11), TO_UNSIGNED( 924, 11), 
		TO_UNSIGNED(1441, 11), TO_UNSIGNED(1477, 11), TO_UNSIGNED( 200, 11), TO_UNSIGNED( 248, 11), TO_UNSIGNED( 817, 11), TO_UNSIGNED( 927, 11), TO_UNSIGNED(1444, 11), TO_UNSIGNED(1465, 11), 
		TO_UNSIGNED( 202, 11), TO_UNSIGNED( 250, 11), TO_UNSIGNED( 823, 11), TO_UNSIGNED( 930, 11), TO_UNSIGNED(1447, 11), TO_UNSIGNED(1471, 11), TO_UNSIGNED( 204, 11), TO_UNSIGNED( 252, 11), 
		TO_UNSIGNED( 829, 11), TO_UNSIGNED( 933, 11), TO_UNSIGNED(1450, 11), TO_UNSIGNED(1495, 11), TO_UNSIGNED( 206, 11), TO_UNSIGNED( 254, 11), TO_UNSIGNED( 691, 11), TO_UNSIGNED( 936, 11), 
		TO_UNSIGNED(1453, 11), TO_UNSIGNED(1501, 11), TO_UNSIGNED( 208, 11), TO_UNSIGNED( 256, 11), TO_UNSIGNED( 697, 11), TO_UNSIGNED( 939, 11), TO_UNSIGNED(1456, 11), TO_UNSIGNED(1507, 11), 
		TO_UNSIGNED( 210, 11), TO_UNSIGNED( 258, 11), TO_UNSIGNED( 703, 11), TO_UNSIGNED( 942, 11), TO_UNSIGNED(1462, 11), TO_UNSIGNED(1489, 11), TO_UNSIGNED( 212, 11), TO_UNSIGNED( 260, 11), 
		TO_UNSIGNED( 709, 11), TO_UNSIGNED( 945, 11), TO_UNSIGNED(1459, 11), TO_UNSIGNED(1513, 11), TO_UNSIGNED( 214, 11), TO_UNSIGNED( 262, 11), TO_UNSIGNED( 715, 11), TO_UNSIGNED( 948, 11), 
		TO_UNSIGNED(1486, 11), TO_UNSIGNED(1525, 11), TO_UNSIGNED( 216, 11), TO_UNSIGNED( 264, 11), TO_UNSIGNED( 721, 11), TO_UNSIGNED( 951, 11), TO_UNSIGNED(1519, 11), TO_UNSIGNED(1618, 11), 
		TO_UNSIGNED( 218, 11), TO_UNSIGNED( 266, 11), TO_UNSIGNED( 727, 11), TO_UNSIGNED( 954, 11), TO_UNSIGNED(1399, 11), TO_UNSIGNED(1543, 11), TO_UNSIGNED( 220, 11), TO_UNSIGNED( 268, 11), 
		TO_UNSIGNED( 733, 11), TO_UNSIGNED( 957, 11), TO_UNSIGNED(1402, 11), TO_UNSIGNED(1549, 11), TO_UNSIGNED( 222, 11), TO_UNSIGNED( 270, 11), TO_UNSIGNED( 739, 11), TO_UNSIGNED( 960, 11), 
		TO_UNSIGNED(1405, 11), TO_UNSIGNED(1531, 11), TO_UNSIGNED( 224, 11), TO_UNSIGNED( 272, 11), TO_UNSIGNED( 745, 11), TO_UNSIGNED( 963, 11), TO_UNSIGNED(1414, 11), TO_UNSIGNED(1537, 11), 
		TO_UNSIGNED( 226, 11), TO_UNSIGNED( 274, 11), TO_UNSIGNED( 751, 11), TO_UNSIGNED( 966, 11), TO_UNSIGNED(1417, 11), TO_UNSIGNED(1555, 11), TO_UNSIGNED( 228, 11), TO_UNSIGNED( 276, 11), 
		TO_UNSIGNED( 757, 11), TO_UNSIGNED( 969, 11), TO_UNSIGNED(1420, 11), TO_UNSIGNED(1561, 11), TO_UNSIGNED( 230, 11), TO_UNSIGNED( 278, 11), TO_UNSIGNED( 763, 11), TO_UNSIGNED( 972, 11), 
		TO_UNSIGNED(1408, 11), TO_UNSIGNED(1573, 11), TO_UNSIGNED( 232, 11), TO_UNSIGNED( 280, 11), TO_UNSIGNED( 769, 11), TO_UNSIGNED( 975, 11), TO_UNSIGNED(1411, 11), TO_UNSIGNED(1567, 11), 
		TO_UNSIGNED( 235, 11), TO_UNSIGNED( 282, 11), TO_UNSIGNED( 788, 11), TO_UNSIGNED(1206, 11), TO_UNSIGNED(1556, 11), TO_UNSIGNED(1635, 11), TO_UNSIGNED( 237, 11), TO_UNSIGNED( 284, 11), 
		TO_UNSIGNED( 794, 11), TO_UNSIGNED(1209, 11), TO_UNSIGNED(1562, 11), TO_UNSIGNED(1629, 11), TO_UNSIGNED( 239, 11), TO_UNSIGNED( 286, 11), TO_UNSIGNED( 800, 11), TO_UNSIGNED(1194, 11), 
		TO_UNSIGNED(1574, 11), TO_UNSIGNED(1632, 11), TO_UNSIGNED( 241, 11), TO_UNSIGNED( 288, 11), TO_UNSIGNED( 806, 11), TO_UNSIGNED(1215, 11), TO_UNSIGNED(1568, 11), TO_UNSIGNED(1641, 11), 
		TO_UNSIGNED( 243, 11), TO_UNSIGNED( 290, 11), TO_UNSIGNED( 812, 11), TO_UNSIGNED(1212, 11), TO_UNSIGNED(1586, 11), TO_UNSIGNED(1638, 11), TO_UNSIGNED( 245, 11), TO_UNSIGNED( 292, 11), 
		TO_UNSIGNED( 818, 11), TO_UNSIGNED(1221, 11), TO_UNSIGNED(1580, 11), TO_UNSIGNED(1644, 11), TO_UNSIGNED( 247, 11), TO_UNSIGNED( 294, 11), TO_UNSIGNED( 824, 11), TO_UNSIGNED(1224, 11), 
		TO_UNSIGNED(1598, 11), TO_UNSIGNED(1650, 11), TO_UNSIGNED( 249, 11), TO_UNSIGNED( 296, 11), TO_UNSIGNED( 830, 11), TO_UNSIGNED(1227, 11), TO_UNSIGNED(1604, 11), TO_UNSIGNED(1647, 11), 
		TO_UNSIGNED( 251, 11), TO_UNSIGNED( 298, 11), TO_UNSIGNED( 692, 11), TO_UNSIGNED(1218, 11), TO_UNSIGNED(1592, 11), TO_UNSIGNED(1653, 11), TO_UNSIGNED(   2, 11), TO_UNSIGNED( 253, 11), 
		TO_UNSIGNED( 300, 11), TO_UNSIGNED( 698, 11), TO_UNSIGNED(1233, 11), TO_UNSIGNED(1656, 11), TO_UNSIGNED( 255, 11), TO_UNSIGNED( 302, 11), TO_UNSIGNED( 704, 11), TO_UNSIGNED(1236, 11), 
		TO_UNSIGNED(1478, 11), TO_UNSIGNED(1659, 11), TO_UNSIGNED( 257, 11), TO_UNSIGNED( 304, 11), TO_UNSIGNED( 710, 11), TO_UNSIGNED(1239, 11), TO_UNSIGNED(1466, 11), TO_UNSIGNED(1662, 11), 
		TO_UNSIGNED( 259, 11), TO_UNSIGNED( 306, 11), TO_UNSIGNED( 716, 11), TO_UNSIGNED(1230, 11), TO_UNSIGNED(1472, 11), TO_UNSIGNED(1665, 11), TO_UNSIGNED( 261, 11), TO_UNSIGNED( 308, 11), 
		TO_UNSIGNED( 722, 11), TO_UNSIGNED(1251, 11), TO_UNSIGNED(1496, 11), TO_UNSIGNED(1671, 11), TO_UNSIGNED( 263, 11), TO_UNSIGNED( 310, 11), TO_UNSIGNED( 728, 11), TO_UNSIGNED(1242, 11), 
		TO_UNSIGNED(1502, 11), TO_UNSIGNED(1668, 11), TO_UNSIGNED( 265, 11), TO_UNSIGNED( 312, 11), TO_UNSIGNED( 734, 11), TO_UNSIGNED(1245, 11), TO_UNSIGNED(1508, 11), TO_UNSIGNED(1674, 11), 
		TO_UNSIGNED( 267, 11), TO_UNSIGNED( 314, 11), TO_UNSIGNED( 740, 11), TO_UNSIGNED(1248, 11), TO_UNSIGNED(1490, 11), TO_UNSIGNED(1677, 11), TO_UNSIGNED( 269, 11), TO_UNSIGNED( 316, 11), 
		TO_UNSIGNED( 746, 11), TO_UNSIGNED(1257, 11), TO_UNSIGNED(1514, 11), TO_UNSIGNED(1680, 11), TO_UNSIGNED( 271, 11), TO_UNSIGNED( 318, 11), TO_UNSIGNED( 752, 11), TO_UNSIGNED(1254, 11), 
		TO_UNSIGNED(1482, 11), TO_UNSIGNED(1526, 11), TO_UNSIGNED( 273, 11), TO_UNSIGNED( 320, 11), TO_UNSIGNED( 758, 11), TO_UNSIGNED(1263, 11), TO_UNSIGNED(1520, 11), TO_UNSIGNED(1608, 11), 
		TO_UNSIGNED( 275, 11), TO_UNSIGNED( 322, 11), TO_UNSIGNED( 764, 11), TO_UNSIGNED(1260, 11), TO_UNSIGNED(1544, 11), TO_UNSIGNED(1611, 11), TO_UNSIGNED( 277, 11), TO_UNSIGNED( 324, 11), 
		TO_UNSIGNED( 770, 11), TO_UNSIGNED(1197, 11), TO_UNSIGNED(1550, 11), TO_UNSIGNED(1620, 11), TO_UNSIGNED( 279, 11), TO_UNSIGNED( 326, 11), TO_UNSIGNED( 776, 11), TO_UNSIGNED(1200, 11), 
		TO_UNSIGNED(1532, 11), TO_UNSIGNED(1623, 11), TO_UNSIGNED( 281, 11), TO_UNSIGNED( 328, 11), TO_UNSIGNED( 782, 11), TO_UNSIGNED(1203, 11), TO_UNSIGNED(1538, 11), TO_UNSIGNED(1626, 11), 
		TO_UNSIGNED( 330, 11), TO_UNSIGNED( 378, 11), TO_UNSIGNED( 705, 11), TO_UNSIGNED( 885, 11), TO_UNSIGNED(1605, 11), TO_UNSIGNED(1669, 11), TO_UNSIGNED( 332, 11), TO_UNSIGNED( 380, 11), 
		TO_UNSIGNED( 711, 11), TO_UNSIGNED( 888, 11), TO_UNSIGNED(1593, 11), TO_UNSIGNED(1675, 11), TO_UNSIGNED(   3, 11), TO_UNSIGNED( 334, 11), TO_UNSIGNED( 382, 11), TO_UNSIGNED( 717, 11), 
		TO_UNSIGNED( 891, 11), TO_UNSIGNED(1678, 11), TO_UNSIGNED( 336, 11), TO_UNSIGNED( 384, 11), TO_UNSIGNED( 723, 11), TO_UNSIGNED( 894, 11), TO_UNSIGNED(1479, 11), TO_UNSIGNED(1681, 11), 
		TO_UNSIGNED( 338, 11), TO_UNSIGNED( 386, 11), TO_UNSIGNED( 729, 11), TO_UNSIGNED( 897, 11), TO_UNSIGNED(1467, 11), TO_UNSIGNED(1483, 11), TO_UNSIGNED( 340, 11), TO_UNSIGNED( 388, 11), 
		TO_UNSIGNED( 735, 11), TO_UNSIGNED( 900, 11), TO_UNSIGNED(1473, 11), TO_UNSIGNED(1609, 11), TO_UNSIGNED( 342, 11), TO_UNSIGNED( 390, 11), TO_UNSIGNED( 741, 11), TO_UNSIGNED( 903, 11), 
		TO_UNSIGNED(1497, 11), TO_UNSIGNED(1612, 11), TO_UNSIGNED( 344, 11), TO_UNSIGNED( 392, 11), TO_UNSIGNED( 747, 11), TO_UNSIGNED( 834, 11), TO_UNSIGNED(1503, 11), TO_UNSIGNED(1621, 11), 
		TO_UNSIGNED( 346, 11), TO_UNSIGNED( 394, 11), TO_UNSIGNED( 753, 11), TO_UNSIGNED( 837, 11), TO_UNSIGNED(1509, 11), TO_UNSIGNED(1624, 11), TO_UNSIGNED( 348, 11), TO_UNSIGNED( 396, 11), 
		TO_UNSIGNED( 759, 11), TO_UNSIGNED( 840, 11), TO_UNSIGNED(1491, 11), TO_UNSIGNED(1627, 11), TO_UNSIGNED( 350, 11), TO_UNSIGNED( 398, 11), TO_UNSIGNED( 765, 11), TO_UNSIGNED( 843, 11), 
		TO_UNSIGNED(1515, 11), TO_UNSIGNED(1636, 11), TO_UNSIGNED( 352, 11), TO_UNSIGNED( 400, 11), TO_UNSIGNED( 771, 11), TO_UNSIGNED( 846, 11), TO_UNSIGNED(1527, 11), TO_UNSIGNED(1630, 11), 
		TO_UNSIGNED( 354, 11), TO_UNSIGNED( 402, 11), TO_UNSIGNED( 777, 11), TO_UNSIGNED( 849, 11), TO_UNSIGNED(1521, 11), TO_UNSIGNED(1633, 11), TO_UNSIGNED( 356, 11), TO_UNSIGNED( 404, 11), 
		TO_UNSIGNED( 783, 11), TO_UNSIGNED( 852, 11), TO_UNSIGNED(1545, 11), TO_UNSIGNED(1642, 11), TO_UNSIGNED( 358, 11), TO_UNSIGNED( 406, 11), TO_UNSIGNED( 789, 11), TO_UNSIGNED( 855, 11), 
		TO_UNSIGNED(1551, 11), TO_UNSIGNED(1639, 11), TO_UNSIGNED( 360, 11), TO_UNSIGNED( 408, 11), TO_UNSIGNED( 795, 11), TO_UNSIGNED( 858, 11), TO_UNSIGNED(1533, 11), TO_UNSIGNED(1645, 11), 
		TO_UNSIGNED( 362, 11), TO_UNSIGNED( 410, 11), TO_UNSIGNED( 801, 11), TO_UNSIGNED( 861, 11), TO_UNSIGNED(1539, 11), TO_UNSIGNED(1651, 11), TO_UNSIGNED( 364, 11), TO_UNSIGNED( 412, 11), 
		TO_UNSIGNED( 807, 11), TO_UNSIGNED( 864, 11), TO_UNSIGNED(1557, 11), TO_UNSIGNED(1648, 11), TO_UNSIGNED( 366, 11), TO_UNSIGNED( 414, 11), TO_UNSIGNED( 813, 11), TO_UNSIGNED( 867, 11), 
		TO_UNSIGNED(1563, 11), TO_UNSIGNED(1654, 11), TO_UNSIGNED( 368, 11), TO_UNSIGNED( 416, 11), TO_UNSIGNED( 819, 11), TO_UNSIGNED( 870, 11), TO_UNSIGNED(1575, 11), TO_UNSIGNED(1657, 11), 
		TO_UNSIGNED( 370, 11), TO_UNSIGNED( 418, 11), TO_UNSIGNED( 825, 11), TO_UNSIGNED( 873, 11), TO_UNSIGNED(1569, 11), TO_UNSIGNED(1660, 11), TO_UNSIGNED( 372, 11), TO_UNSIGNED( 420, 11), 
		TO_UNSIGNED( 831, 11), TO_UNSIGNED( 876, 11), TO_UNSIGNED(1587, 11), TO_UNSIGNED(1663, 11), TO_UNSIGNED( 374, 11), TO_UNSIGNED( 422, 11), TO_UNSIGNED( 693, 11), TO_UNSIGNED( 879, 11), 
		TO_UNSIGNED(1581, 11), TO_UNSIGNED(1666, 11), TO_UNSIGNED( 376, 11), TO_UNSIGNED( 424, 11), TO_UNSIGNED( 699, 11), TO_UNSIGNED( 882, 11), TO_UNSIGNED(1599, 11), TO_UNSIGNED(1672, 11), 
		TO_UNSIGNED( 379, 11), TO_UNSIGNED( 426, 11), TO_UNSIGNED( 682, 11), TO_UNSIGNED( 736, 11), TO_UNSIGNED(1198, 11), TO_UNSIGNED(1540, 11), TO_UNSIGNED( 381, 11), TO_UNSIGNED( 428, 11), 
		TO_UNSIGNED( 685, 11), TO_UNSIGNED( 742, 11), TO_UNSIGNED(1201, 11), TO_UNSIGNED(1558, 11), TO_UNSIGNED( 383, 11), TO_UNSIGNED( 430, 11), TO_UNSIGNED( 688, 11), TO_UNSIGNED( 748, 11), 
		TO_UNSIGNED(1204, 11), TO_UNSIGNED(1564, 11), TO_UNSIGNED( 385, 11), TO_UNSIGNED( 432, 11), TO_UNSIGNED( 619, 11), TO_UNSIGNED( 754, 11), TO_UNSIGNED(1207, 11), TO_UNSIGNED(1576, 11), 
		TO_UNSIGNED( 387, 11), TO_UNSIGNED( 434, 11), TO_UNSIGNED( 622, 11), TO_UNSIGNED( 760, 11), TO_UNSIGNED(1210, 11), TO_UNSIGNED(1570, 11), TO_UNSIGNED( 389, 11), TO_UNSIGNED( 436, 11), 
		TO_UNSIGNED( 625, 11), TO_UNSIGNED( 766, 11), TO_UNSIGNED(1195, 11), TO_UNSIGNED(1588, 11), TO_UNSIGNED( 391, 11), TO_UNSIGNED( 438, 11), TO_UNSIGNED( 628, 11), TO_UNSIGNED( 772, 11), 
		TO_UNSIGNED(1216, 11), TO_UNSIGNED(1582, 11), TO_UNSIGNED( 393, 11), TO_UNSIGNED( 440, 11), TO_UNSIGNED( 631, 11), TO_UNSIGNED( 778, 11), TO_UNSIGNED(1213, 11), TO_UNSIGNED(1600, 11), 
		TO_UNSIGNED( 395, 11), TO_UNSIGNED( 442, 11), TO_UNSIGNED( 634, 11), TO_UNSIGNED( 784, 11), TO_UNSIGNED(1222, 11), TO_UNSIGNED(1606, 11), TO_UNSIGNED( 397, 11), TO_UNSIGNED( 444, 11), 
		TO_UNSIGNED( 637, 11), TO_UNSIGNED( 790, 11), TO_UNSIGNED(1225, 11), TO_UNSIGNED(1594, 11), TO_UNSIGNED(   4, 11), TO_UNSIGNED( 399, 11), TO_UNSIGNED( 446, 11), TO_UNSIGNED( 640, 11), 
		TO_UNSIGNED( 796, 11), TO_UNSIGNED(1228, 11), TO_UNSIGNED( 401, 11), TO_UNSIGNED( 448, 11), TO_UNSIGNED( 643, 11), TO_UNSIGNED( 802, 11), TO_UNSIGNED(1219, 11), TO_UNSIGNED(1480, 11), 
		TO_UNSIGNED( 403, 11), TO_UNSIGNED( 450, 11), TO_UNSIGNED( 646, 11), TO_UNSIGNED( 808, 11), TO_UNSIGNED(1234, 11), TO_UNSIGNED(1468, 11), TO_UNSIGNED( 405, 11), TO_UNSIGNED( 452, 11), 
		TO_UNSIGNED( 649, 11), TO_UNSIGNED( 814, 11), TO_UNSIGNED(1237, 11), TO_UNSIGNED(1474, 11), TO_UNSIGNED( 407, 11), TO_UNSIGNED( 454, 11), TO_UNSIGNED( 652, 11), TO_UNSIGNED( 820, 11), 
		TO_UNSIGNED(1240, 11), TO_UNSIGNED(1498, 11), TO_UNSIGNED( 409, 11), TO_UNSIGNED( 456, 11), TO_UNSIGNED( 655, 11), TO_UNSIGNED( 826, 11), TO_UNSIGNED(1231, 11), TO_UNSIGNED(1504, 11), 
		TO_UNSIGNED( 411, 11), TO_UNSIGNED( 458, 11), TO_UNSIGNED( 658, 11), TO_UNSIGNED( 832, 11), TO_UNSIGNED(1252, 11), TO_UNSIGNED(1510, 11), TO_UNSIGNED( 413, 11), TO_UNSIGNED( 460, 11), 
		TO_UNSIGNED( 661, 11), TO_UNSIGNED( 694, 11), TO_UNSIGNED(1243, 11), TO_UNSIGNED(1492, 11), TO_UNSIGNED( 415, 11), TO_UNSIGNED( 462, 11), TO_UNSIGNED( 664, 11), TO_UNSIGNED( 700, 11), 
		TO_UNSIGNED(1246, 11), TO_UNSIGNED(1516, 11), TO_UNSIGNED( 417, 11), TO_UNSIGNED( 464, 11), TO_UNSIGNED( 667, 11), TO_UNSIGNED( 706, 11), TO_UNSIGNED(1249, 11), TO_UNSIGNED(1528, 11), 
		TO_UNSIGNED( 419, 11), TO_UNSIGNED( 466, 11), TO_UNSIGNED( 670, 11), TO_UNSIGNED( 712, 11), TO_UNSIGNED(1258, 11), TO_UNSIGNED(1522, 11), TO_UNSIGNED( 421, 11), TO_UNSIGNED( 468, 11), 
		TO_UNSIGNED( 673, 11), TO_UNSIGNED( 718, 11), TO_UNSIGNED(1255, 11), TO_UNSIGNED(1546, 11), TO_UNSIGNED( 423, 11), TO_UNSIGNED( 470, 11), TO_UNSIGNED( 676, 11), TO_UNSIGNED( 724, 11), 
		TO_UNSIGNED(1264, 11), TO_UNSIGNED(1552, 11), TO_UNSIGNED( 425, 11), TO_UNSIGNED( 472, 11), TO_UNSIGNED( 679, 11), TO_UNSIGNED( 730, 11), TO_UNSIGNED(1261, 11), TO_UNSIGNED(1534, 11), 
		TO_UNSIGNED( 474, 11), TO_UNSIGNED( 522, 11), TO_UNSIGNED(1062, 11), TO_UNSIGNED(1332, 11), TO_UNSIGNED(1631, 11), TO_UNSIGNED(1729, 11), TO_UNSIGNED( 476, 11), TO_UNSIGNED( 524, 11), 
		TO_UNSIGNED(1068, 11), TO_UNSIGNED(1326, 11), TO_UNSIGNED(1634, 11), TO_UNSIGNED(1723, 11), TO_UNSIGNED( 478, 11), TO_UNSIGNED( 526, 11), TO_UNSIGNED(1074, 11), TO_UNSIGNED(1350, 11), 
		TO_UNSIGNED(1643, 11), TO_UNSIGNED(1735, 11), TO_UNSIGNED( 480, 11), TO_UNSIGNED( 528, 11), TO_UNSIGNED(1080, 11), TO_UNSIGNED(1356, 11), TO_UNSIGNED(1640, 11), TO_UNSIGNED(1771, 11), 
		TO_UNSIGNED( 482, 11), TO_UNSIGNED( 530, 11), TO_UNSIGNED(1086, 11), TO_UNSIGNED(1338, 11), TO_UNSIGNED(1646, 11), TO_UNSIGNED(1777, 11), TO_UNSIGNED( 484, 11), TO_UNSIGNED( 532, 11), 
		TO_UNSIGNED(1092, 11), TO_UNSIGNED(1344, 11), TO_UNSIGNED(1652, 11), TO_UNSIGNED(1741, 11), TO_UNSIGNED( 486, 11), TO_UNSIGNED( 534, 11), TO_UNSIGNED(1098, 11), TO_UNSIGNED(1368, 11), 
		TO_UNSIGNED(1649, 11), TO_UNSIGNED(1747, 11), TO_UNSIGNED( 488, 11), TO_UNSIGNED( 536, 11), TO_UNSIGNED(1104, 11), TO_UNSIGNED(1374, 11), TO_UNSIGNED(1655, 11), TO_UNSIGNED(1753, 11), 
		TO_UNSIGNED( 490, 11), TO_UNSIGNED( 538, 11), TO_UNSIGNED(1110, 11), TO_UNSIGNED(1362, 11), TO_UNSIGNED(1658, 11), TO_UNSIGNED(1759, 11), TO_UNSIGNED( 492, 11), TO_UNSIGNED( 540, 11), 
		TO_UNSIGNED(1116, 11), TO_UNSIGNED(1392, 11), TO_UNSIGNED(1661, 11), TO_UNSIGNED(1765, 11), TO_UNSIGNED( 494, 11), TO_UNSIGNED( 542, 11), TO_UNSIGNED( 978, 11), TO_UNSIGNED(1380, 11), 
		TO_UNSIGNED(1664, 11), TO_UNSIGNED(1801, 11), TO_UNSIGNED( 496, 11), TO_UNSIGNED( 544, 11), TO_UNSIGNED( 984, 11), TO_UNSIGNED(1386, 11), TO_UNSIGNED(1667, 11), TO_UNSIGNED(1789, 11), 
		TO_UNSIGNED( 130, 11), TO_UNSIGNED( 498, 11), TO_UNSIGNED( 546, 11), TO_UNSIGNED( 990, 11), TO_UNSIGNED(1673, 11), TO_UNSIGNED(1795, 11), TO_UNSIGNED(  78, 11), TO_UNSIGNED( 500, 11), 
		TO_UNSIGNED( 548, 11), TO_UNSIGNED( 996, 11), TO_UNSIGNED(1670, 11), TO_UNSIGNED(1807, 11), TO_UNSIGNED( 502, 11), TO_UNSIGNED( 550, 11), TO_UNSIGNED(1002, 11), TO_UNSIGNED(1272, 11), 
		TO_UNSIGNED(1676, 11), TO_UNSIGNED(1783, 11), TO_UNSIGNED(   6, 11), TO_UNSIGNED( 504, 11), TO_UNSIGNED( 552, 11), TO_UNSIGNED(1008, 11), TO_UNSIGNED(1278, 11), TO_UNSIGNED(1679, 11), 
		TO_UNSIGNED( 506, 11), TO_UNSIGNED( 554, 11), TO_UNSIGNED(1014, 11), TO_UNSIGNED(1284, 11), TO_UNSIGNED(1682, 11), TO_UNSIGNED(1813, 11), TO_UNSIGNED( 136, 11), TO_UNSIGNED( 508, 11), 
		TO_UNSIGNED( 556, 11), TO_UNSIGNED(1020, 11), TO_UNSIGNED(1266, 11), TO_UNSIGNED(1484, 11), TO_UNSIGNED( 510, 11), TO_UNSIGNED( 558, 11), TO_UNSIGNED(1026, 11), TO_UNSIGNED(1296, 11), 
		TO_UNSIGNED(1610, 11), TO_UNSIGNED(1687, 11), TO_UNSIGNED( 512, 11), TO_UNSIGNED( 560, 11), TO_UNSIGNED(1032, 11), TO_UNSIGNED(1290, 11), TO_UNSIGNED(1613, 11), TO_UNSIGNED(1711, 11), 
		TO_UNSIGNED( 514, 11), TO_UNSIGNED( 562, 11), TO_UNSIGNED(1038, 11), TO_UNSIGNED(1308, 11), TO_UNSIGNED(1622, 11), TO_UNSIGNED(1699, 11), TO_UNSIGNED( 516, 11), TO_UNSIGNED( 564, 11), 
		TO_UNSIGNED(1044, 11), TO_UNSIGNED(1302, 11), TO_UNSIGNED(1625, 11), TO_UNSIGNED(1705, 11), TO_UNSIGNED( 518, 11), TO_UNSIGNED( 566, 11), TO_UNSIGNED(1050, 11), TO_UNSIGNED(1314, 11), 
		TO_UNSIGNED(1628, 11), TO_UNSIGNED(1693, 11), TO_UNSIGNED( 520, 11), TO_UNSIGNED( 568, 11), TO_UNSIGNED(1056, 11), TO_UNSIGNED(1320, 11), TO_UNSIGNED(1637, 11), TO_UNSIGNED(1717, 11), 
		TO_UNSIGNED( 523, 11), TO_UNSIGNED( 570, 11), TO_UNSIGNED( 695, 11), TO_UNSIGNED( 877, 11), TO_UNSIGNED(1445, 11), TO_UNSIGNED(1535, 11), TO_UNSIGNED( 525, 11), TO_UNSIGNED( 572, 11), 
		TO_UNSIGNED( 701, 11), TO_UNSIGNED( 880, 11), TO_UNSIGNED(1448, 11), TO_UNSIGNED(1541, 11), TO_UNSIGNED( 527, 11), TO_UNSIGNED( 574, 11), TO_UNSIGNED( 707, 11), TO_UNSIGNED( 883, 11), 
		TO_UNSIGNED(1451, 11), TO_UNSIGNED(1559, 11), TO_UNSIGNED( 529, 11), TO_UNSIGNED( 576, 11), TO_UNSIGNED( 713, 11), TO_UNSIGNED( 886, 11), TO_UNSIGNED(1454, 11), TO_UNSIGNED(1565, 11), 
		TO_UNSIGNED( 531, 11), TO_UNSIGNED( 578, 11), TO_UNSIGNED( 719, 11), TO_UNSIGNED( 889, 11), TO_UNSIGNED(1457, 11), TO_UNSIGNED(1577, 11), TO_UNSIGNED( 533, 11), TO_UNSIGNED( 580, 11), 
		TO_UNSIGNED( 725, 11), TO_UNSIGNED( 892, 11), TO_UNSIGNED(1463, 11), TO_UNSIGNED(1571, 11), TO_UNSIGNED( 535, 11), TO_UNSIGNED( 582, 11), TO_UNSIGNED( 731, 11), TO_UNSIGNED( 895, 11), 
		TO_UNSIGNED(1460, 11), TO_UNSIGNED(1589, 11), TO_UNSIGNED( 537, 11), TO_UNSIGNED( 584, 11), TO_UNSIGNED( 737, 11), TO_UNSIGNED( 898, 11), TO_UNSIGNED(1487, 11), TO_UNSIGNED(1583, 11), 
		TO_UNSIGNED( 539, 11), TO_UNSIGNED( 586, 11), TO_UNSIGNED( 743, 11), TO_UNSIGNED( 901, 11), TO_UNSIGNED(1601, 11), TO_UNSIGNED(1619, 11), TO_UNSIGNED( 541, 11), TO_UNSIGNED( 588, 11), 
		TO_UNSIGNED( 749, 11), TO_UNSIGNED( 904, 11), TO_UNSIGNED(1400, 11), TO_UNSIGNED(1607, 11), TO_UNSIGNED( 543, 11), TO_UNSIGNED( 590, 11), TO_UNSIGNED( 755, 11), TO_UNSIGNED( 835, 11), 
		TO_UNSIGNED(1403, 11), TO_UNSIGNED(1595, 11), TO_UNSIGNED(   5, 11), TO_UNSIGNED( 545, 11), TO_UNSIGNED( 592, 11), TO_UNSIGNED( 761, 11), TO_UNSIGNED( 838, 11), TO_UNSIGNED(1406, 11), 
		TO_UNSIGNED( 547, 11), TO_UNSIGNED( 594, 11), TO_UNSIGNED( 767, 11), TO_UNSIGNED( 841, 11), TO_UNSIGNED(1415, 11), TO_UNSIGNED(1481, 11), TO_UNSIGNED( 549, 11), TO_UNSIGNED( 596, 11), 
		TO_UNSIGNED( 773, 11), TO_UNSIGNED( 844, 11), TO_UNSIGNED(1418, 11), TO_UNSIGNED(1469, 11), TO_UNSIGNED( 551, 11), TO_UNSIGNED( 598, 11), TO_UNSIGNED( 779, 11), TO_UNSIGNED( 847, 11), 
		TO_UNSIGNED(1421, 11), TO_UNSIGNED(1475, 11), TO_UNSIGNED( 553, 11), TO_UNSIGNED( 600, 11), TO_UNSIGNED( 785, 11), TO_UNSIGNED( 850, 11), TO_UNSIGNED(1409, 11), TO_UNSIGNED(1499, 11), 
		TO_UNSIGNED( 555, 11), TO_UNSIGNED( 602, 11), TO_UNSIGNED( 791, 11), TO_UNSIGNED( 853, 11), TO_UNSIGNED(1412, 11), TO_UNSIGNED(1505, 11), TO_UNSIGNED( 557, 11), TO_UNSIGNED( 604, 11), 
		TO_UNSIGNED( 797, 11), TO_UNSIGNED( 856, 11), TO_UNSIGNED(1436, 11), TO_UNSIGNED(1511, 11), TO_UNSIGNED( 559, 11), TO_UNSIGNED( 606, 11), TO_UNSIGNED( 803, 11), TO_UNSIGNED( 859, 11), 
		TO_UNSIGNED(1433, 11), TO_UNSIGNED(1493, 11), TO_UNSIGNED( 561, 11), TO_UNSIGNED( 608, 11), TO_UNSIGNED( 809, 11), TO_UNSIGNED( 862, 11), TO_UNSIGNED(1424, 11), TO_UNSIGNED(1517, 11), 
		TO_UNSIGNED( 563, 11), TO_UNSIGNED( 610, 11), TO_UNSIGNED( 815, 11), TO_UNSIGNED( 865, 11), TO_UNSIGNED(1427, 11), TO_UNSIGNED(1529, 11), TO_UNSIGNED( 565, 11), TO_UNSIGNED( 612, 11), 
		TO_UNSIGNED( 821, 11), TO_UNSIGNED( 868, 11), TO_UNSIGNED(1430, 11), TO_UNSIGNED(1523, 11), TO_UNSIGNED( 567, 11), TO_UNSIGNED( 614, 11), TO_UNSIGNED( 827, 11), TO_UNSIGNED( 871, 11), 
		TO_UNSIGNED(1439, 11), TO_UNSIGNED(1547, 11), TO_UNSIGNED( 569, 11), TO_UNSIGNED( 616, 11), TO_UNSIGNED( 833, 11), TO_UNSIGNED( 874, 11), TO_UNSIGNED(1442, 11), TO_UNSIGNED(1553, 11), 
		TO_UNSIGNED(  76, 11), TO_UNSIGNED( 571, 11), TO_UNSIGNED( 922, 11), TO_UNSIGNED(1105, 11), TO_UNSIGNED(1339, 11), TO_UNSIGNED(1796, 11), TO_UNSIGNED( 573, 11), TO_UNSIGNED( 925, 11), 
		TO_UNSIGNED(1111, 11), TO_UNSIGNED(1345, 11), TO_UNSIGNED(1615, 11), TO_UNSIGNED(1808, 11), TO_UNSIGNED( 575, 11), TO_UNSIGNED( 928, 11), TO_UNSIGNED(1117, 11), TO_UNSIGNED(1369, 11), 
		TO_UNSIGNED(1784, 11), TO_UNSIGNED(1820, 11), TO_UNSIGNED(   7, 11), TO_UNSIGNED(  13, 11), TO_UNSIGNED( 577, 11), TO_UNSIGNED( 931, 11), TO_UNSIGNED( 979, 11), TO_UNSIGNED(1375, 11), 
		TO_UNSIGNED(  16, 11), TO_UNSIGNED( 579, 11), TO_UNSIGNED( 934, 11), TO_UNSIGNED( 985, 11), TO_UNSIGNED(1363, 11), TO_UNSIGNED(1814, 11), TO_UNSIGNED(  19, 11), TO_UNSIGNED( 137, 11), 
		TO_UNSIGNED( 581, 11), TO_UNSIGNED( 937, 11), TO_UNSIGNED( 991, 11), TO_UNSIGNED(1393, 11), TO_UNSIGNED(  22, 11), TO_UNSIGNED( 583, 11), TO_UNSIGNED( 940, 11), TO_UNSIGNED( 997, 11), 
		TO_UNSIGNED(1381, 11), TO_UNSIGNED(1688, 11), TO_UNSIGNED(  25, 11), TO_UNSIGNED( 585, 11), TO_UNSIGNED( 943, 11), TO_UNSIGNED(1003, 11), TO_UNSIGNED(1387, 11), TO_UNSIGNED(1712, 11), 
		TO_UNSIGNED(  28, 11), TO_UNSIGNED( 131, 11), TO_UNSIGNED( 587, 11), TO_UNSIGNED( 946, 11), TO_UNSIGNED(1009, 11), TO_UNSIGNED(1700, 11), TO_UNSIGNED(  31, 11), TO_UNSIGNED(  79, 11), 
		TO_UNSIGNED( 589, 11), TO_UNSIGNED( 949, 11), TO_UNSIGNED(1015, 11), TO_UNSIGNED(1706, 11), TO_UNSIGNED(  34, 11), TO_UNSIGNED( 591, 11), TO_UNSIGNED( 952, 11), TO_UNSIGNED(1021, 11), 
		TO_UNSIGNED(1273, 11), TO_UNSIGNED(1694, 11), TO_UNSIGNED(  37, 11), TO_UNSIGNED( 593, 11), TO_UNSIGNED( 955, 11), TO_UNSIGNED(1027, 11), TO_UNSIGNED(1279, 11), TO_UNSIGNED(1718, 11), 
		TO_UNSIGNED(  40, 11), TO_UNSIGNED( 595, 11), TO_UNSIGNED( 958, 11), TO_UNSIGNED(1033, 11), TO_UNSIGNED(1285, 11), TO_UNSIGNED(1730, 11), TO_UNSIGNED(  43, 11), TO_UNSIGNED( 597, 11), 
		TO_UNSIGNED( 961, 11), TO_UNSIGNED(1039, 11), TO_UNSIGNED(1267, 11), TO_UNSIGNED(1724, 11), TO_UNSIGNED(  46, 11), TO_UNSIGNED( 599, 11), TO_UNSIGNED( 964, 11), TO_UNSIGNED(1045, 11), 
		TO_UNSIGNED(1297, 11), TO_UNSIGNED(1736, 11), TO_UNSIGNED(  49, 11), TO_UNSIGNED( 601, 11), TO_UNSIGNED( 967, 11), TO_UNSIGNED(1051, 11), TO_UNSIGNED(1291, 11), TO_UNSIGNED(1772, 11), 
		TO_UNSIGNED(  52, 11), TO_UNSIGNED( 603, 11), TO_UNSIGNED( 970, 11), TO_UNSIGNED(1057, 11), TO_UNSIGNED(1309, 11), TO_UNSIGNED(1778, 11), TO_UNSIGNED(  55, 11), TO_UNSIGNED( 605, 11), 
		TO_UNSIGNED( 973, 11), TO_UNSIGNED(1063, 11), TO_UNSIGNED(1303, 11), TO_UNSIGNED(1742, 11), TO_UNSIGNED(  58, 11), TO_UNSIGNED( 607, 11), TO_UNSIGNED( 976, 11), TO_UNSIGNED(1069, 11), 
		TO_UNSIGNED(1315, 11), TO_UNSIGNED(1748, 11), TO_UNSIGNED(  61, 11), TO_UNSIGNED( 609, 11), TO_UNSIGNED( 907, 11), TO_UNSIGNED(1075, 11), TO_UNSIGNED(1321, 11), TO_UNSIGNED(1754, 11), 
		TO_UNSIGNED(  64, 11), TO_UNSIGNED( 611, 11), TO_UNSIGNED( 910, 11), TO_UNSIGNED(1081, 11), TO_UNSIGNED(1333, 11), TO_UNSIGNED(1760, 11), TO_UNSIGNED(  67, 11), TO_UNSIGNED( 613, 11), 
		TO_UNSIGNED( 913, 11), TO_UNSIGNED(1087, 11), TO_UNSIGNED(1327, 11), TO_UNSIGNED(1766, 11), TO_UNSIGNED(  70, 11), TO_UNSIGNED( 615, 11), TO_UNSIGNED( 916, 11), TO_UNSIGNED(1093, 11), 
		TO_UNSIGNED(1351, 11), TO_UNSIGNED(1802, 11), TO_UNSIGNED(  73, 11), TO_UNSIGNED( 617, 11), TO_UNSIGNED( 919, 11), TO_UNSIGNED(1099, 11), TO_UNSIGNED(1357, 11), TO_UNSIGNED(1790, 11), 
		TO_UNSIGNED(   8, 11), TO_UNSIGNED( 132, 11), TO_UNSIGNED( 671, 11), TO_UNSIGNED(1028, 11), TO_UNSIGNED(1196, 11), TO_UNSIGNED(1684, 11), TO_UNSIGNED(1685, 11), TO_UNSIGNED(  80, 11), 
		TO_UNSIGNED(  85, 11), TO_UNSIGNED( 674, 11), TO_UNSIGNED(1034, 11), TO_UNSIGNED(1217, 11), TO_UNSIGNED(1815, 11), TO_UNSIGNED(1822, 11), TO_UNSIGNED(  87, 11), TO_UNSIGNED( 138, 11), 
		TO_UNSIGNED( 142, 11), TO_UNSIGNED( 677, 11), TO_UNSIGNED(1040, 11), TO_UNSIGNED(1214, 11), TO_UNSIGNED(1274, 11), TO_UNSIGNED(  89, 11), TO_UNSIGNED( 144, 11), TO_UNSIGNED( 680, 11), 
		TO_UNSIGNED(1046, 11), TO_UNSIGNED(1223, 11), TO_UNSIGNED(1280, 11), TO_UNSIGNED(1689, 11), TO_UNSIGNED(  91, 11), TO_UNSIGNED( 146, 11), TO_UNSIGNED( 683, 11), TO_UNSIGNED(1052, 11), 
		TO_UNSIGNED(1226, 11), TO_UNSIGNED(1286, 11), TO_UNSIGNED(1713, 11), TO_UNSIGNED(  93, 11), TO_UNSIGNED( 148, 11), TO_UNSIGNED( 686, 11), TO_UNSIGNED(1058, 11), TO_UNSIGNED(1229, 11), 
		TO_UNSIGNED(1268, 11), TO_UNSIGNED(1701, 11), TO_UNSIGNED(  95, 11), TO_UNSIGNED( 150, 11), TO_UNSIGNED( 689, 11), TO_UNSIGNED(1064, 11), TO_UNSIGNED(1220, 11), TO_UNSIGNED(1298, 11), 
		TO_UNSIGNED(1707, 11), TO_UNSIGNED(  97, 11), TO_UNSIGNED( 152, 11), TO_UNSIGNED( 620, 11), TO_UNSIGNED(1070, 11), TO_UNSIGNED(1235, 11), TO_UNSIGNED(1292, 11), TO_UNSIGNED(1695, 11), 
		TO_UNSIGNED(  99, 11), TO_UNSIGNED( 154, 11), TO_UNSIGNED( 623, 11), TO_UNSIGNED(1076, 11), TO_UNSIGNED(1238, 11), TO_UNSIGNED(1310, 11), TO_UNSIGNED(1719, 11), TO_UNSIGNED( 101, 11), 
		TO_UNSIGNED( 156, 11), TO_UNSIGNED( 626, 11), TO_UNSIGNED(1082, 11), TO_UNSIGNED(1241, 11), TO_UNSIGNED(1304, 11), TO_UNSIGNED(1731, 11), TO_UNSIGNED( 103, 11), TO_UNSIGNED( 158, 11), 
		TO_UNSIGNED( 629, 11), TO_UNSIGNED(1088, 11), TO_UNSIGNED(1232, 11), TO_UNSIGNED(1316, 11), TO_UNSIGNED(1725, 11), TO_UNSIGNED( 105, 11), TO_UNSIGNED( 160, 11), TO_UNSIGNED( 632, 11), 
		TO_UNSIGNED(1094, 11), TO_UNSIGNED(1253, 11), TO_UNSIGNED(1322, 11), TO_UNSIGNED(1737, 11), TO_UNSIGNED( 107, 11), TO_UNSIGNED( 162, 11), TO_UNSIGNED( 635, 11), TO_UNSIGNED(1100, 11), 
		TO_UNSIGNED(1244, 11), TO_UNSIGNED(1334, 11), TO_UNSIGNED(1773, 11), TO_UNSIGNED( 109, 11), TO_UNSIGNED( 164, 11), TO_UNSIGNED( 638, 11), TO_UNSIGNED(1106, 11), TO_UNSIGNED(1247, 11), 
		TO_UNSIGNED(1328, 11), TO_UNSIGNED(1779, 11), TO_UNSIGNED( 111, 11), TO_UNSIGNED( 166, 11), TO_UNSIGNED( 641, 11), TO_UNSIGNED(1112, 11), TO_UNSIGNED(1250, 11), TO_UNSIGNED(1352, 11), 
		TO_UNSIGNED(1743, 11), TO_UNSIGNED( 113, 11), TO_UNSIGNED( 168, 11), TO_UNSIGNED( 644, 11), TO_UNSIGNED(1118, 11), TO_UNSIGNED(1259, 11), TO_UNSIGNED(1358, 11), TO_UNSIGNED(1749, 11), 
		TO_UNSIGNED( 115, 11), TO_UNSIGNED( 170, 11), TO_UNSIGNED( 647, 11), TO_UNSIGNED( 980, 11), TO_UNSIGNED(1256, 11), TO_UNSIGNED(1340, 11), TO_UNSIGNED(1755, 11), TO_UNSIGNED( 117, 11), 
		TO_UNSIGNED( 172, 11), TO_UNSIGNED( 650, 11), TO_UNSIGNED( 986, 11), TO_UNSIGNED(1265, 11), TO_UNSIGNED(1346, 11), TO_UNSIGNED(1761, 11), TO_UNSIGNED( 119, 11), TO_UNSIGNED( 174, 11), 
		TO_UNSIGNED( 653, 11), TO_UNSIGNED( 992, 11), TO_UNSIGNED(1262, 11), TO_UNSIGNED(1370, 11), TO_UNSIGNED(1767, 11), TO_UNSIGNED( 121, 11), TO_UNSIGNED( 176, 11), TO_UNSIGNED( 656, 11), 
		TO_UNSIGNED( 998, 11), TO_UNSIGNED(1199, 11), TO_UNSIGNED(1376, 11), TO_UNSIGNED(1803, 11), TO_UNSIGNED( 123, 11), TO_UNSIGNED( 178, 11), TO_UNSIGNED( 659, 11), TO_UNSIGNED(1004, 11), 
		TO_UNSIGNED(1202, 11), TO_UNSIGNED(1364, 11), TO_UNSIGNED(1791, 11), TO_UNSIGNED( 125, 11), TO_UNSIGNED( 180, 11), TO_UNSIGNED( 662, 11), TO_UNSIGNED(1010, 11), TO_UNSIGNED(1205, 11), 
		TO_UNSIGNED(1394, 11), TO_UNSIGNED(1797, 11), TO_UNSIGNED( 127, 11), TO_UNSIGNED( 182, 11), TO_UNSIGNED( 665, 11), TO_UNSIGNED(1016, 11), TO_UNSIGNED(1208, 11), TO_UNSIGNED(1382, 11), 
		TO_UNSIGNED(1809, 11), TO_UNSIGNED( 129, 11), TO_UNSIGNED( 184, 11), TO_UNSIGNED( 668, 11), TO_UNSIGNED(1022, 11), TO_UNSIGNED(1211, 11), TO_UNSIGNED(1388, 11), TO_UNSIGNED(1785, 11), 
		TO_UNSIGNED( 187, 11), TO_UNSIGNED( 836, 11), TO_UNSIGNED(1083, 11), TO_UNSIGNED(1140, 11), TO_UNSIGNED(1371, 11), TO_UNSIGNED(1686, 11), TO_UNSIGNED(1690, 11), TO_UNSIGNED( 189, 11), 
		TO_UNSIGNED( 839, 11), TO_UNSIGNED(1089, 11), TO_UNSIGNED(1143, 11), TO_UNSIGNED(1377, 11), TO_UNSIGNED(1714, 11), TO_UNSIGNED(1823, 11), TO_UNSIGNED( 143, 11), TO_UNSIGNED( 191, 11), 
		TO_UNSIGNED( 842, 11), TO_UNSIGNED(1095, 11), TO_UNSIGNED(1146, 11), TO_UNSIGNED(1365, 11), TO_UNSIGNED(1702, 11), TO_UNSIGNED( 145, 11), TO_UNSIGNED( 193, 11), TO_UNSIGNED( 845, 11), 
		TO_UNSIGNED(1101, 11), TO_UNSIGNED(1149, 11), TO_UNSIGNED(1395, 11), TO_UNSIGNED(1708, 11), TO_UNSIGNED( 147, 11), TO_UNSIGNED( 195, 11), TO_UNSIGNED( 848, 11), TO_UNSIGNED(1107, 11), 
		TO_UNSIGNED(1152, 11), TO_UNSIGNED(1383, 11), TO_UNSIGNED(1696, 11), TO_UNSIGNED( 149, 11), TO_UNSIGNED( 197, 11), TO_UNSIGNED( 851, 11), TO_UNSIGNED(1113, 11), TO_UNSIGNED(1155, 11), 
		TO_UNSIGNED(1389, 11), TO_UNSIGNED(1720, 11), TO_UNSIGNED( 133, 11), TO_UNSIGNED( 151, 11), TO_UNSIGNED( 199, 11), TO_UNSIGNED( 854, 11), TO_UNSIGNED(1119, 11), TO_UNSIGNED(1158, 11), 
		TO_UNSIGNED(1732, 11), TO_UNSIGNED(  81, 11), TO_UNSIGNED( 153, 11), TO_UNSIGNED( 201, 11), TO_UNSIGNED( 857, 11), TO_UNSIGNED( 981, 11), TO_UNSIGNED(1161, 11), TO_UNSIGNED(1726, 11), 
		TO_UNSIGNED( 155, 11), TO_UNSIGNED( 203, 11), TO_UNSIGNED( 860, 11), TO_UNSIGNED( 987, 11), TO_UNSIGNED(1164, 11), TO_UNSIGNED(1275, 11), TO_UNSIGNED(1738, 11), TO_UNSIGNED( 157, 11), 
		TO_UNSIGNED( 205, 11), TO_UNSIGNED( 863, 11), TO_UNSIGNED( 993, 11), TO_UNSIGNED(1167, 11), TO_UNSIGNED(1281, 11), TO_UNSIGNED(1774, 11), TO_UNSIGNED( 159, 11), TO_UNSIGNED( 207, 11), 
		TO_UNSIGNED( 866, 11), TO_UNSIGNED( 999, 11), TO_UNSIGNED(1170, 11), TO_UNSIGNED(1287, 11), TO_UNSIGNED(1780, 11), TO_UNSIGNED( 161, 11), TO_UNSIGNED( 209, 11), TO_UNSIGNED( 869, 11), 
		TO_UNSIGNED(1005, 11), TO_UNSIGNED(1173, 11), TO_UNSIGNED(1269, 11), TO_UNSIGNED(1744, 11), TO_UNSIGNED( 163, 11), TO_UNSIGNED( 211, 11), TO_UNSIGNED( 872, 11), TO_UNSIGNED(1011, 11), 
		TO_UNSIGNED(1176, 11), TO_UNSIGNED(1299, 11), TO_UNSIGNED(1750, 11), TO_UNSIGNED( 165, 11), TO_UNSIGNED( 213, 11), TO_UNSIGNED( 875, 11), TO_UNSIGNED(1017, 11), TO_UNSIGNED(1179, 11), 
		TO_UNSIGNED(1293, 11), TO_UNSIGNED(1756, 11), TO_UNSIGNED( 167, 11), TO_UNSIGNED( 215, 11), TO_UNSIGNED( 878, 11), TO_UNSIGNED(1023, 11), TO_UNSIGNED(1182, 11), TO_UNSIGNED(1311, 11), 
		TO_UNSIGNED(1762, 11), TO_UNSIGNED( 169, 11), TO_UNSIGNED( 217, 11), TO_UNSIGNED( 881, 11), TO_UNSIGNED(1029, 11), TO_UNSIGNED(1185, 11), TO_UNSIGNED(1305, 11), TO_UNSIGNED(1768, 11), 
		TO_UNSIGNED( 171, 11), TO_UNSIGNED( 219, 11), TO_UNSIGNED( 884, 11), TO_UNSIGNED(1035, 11), TO_UNSIGNED(1188, 11), TO_UNSIGNED(1317, 11), TO_UNSIGNED(1804, 11), TO_UNSIGNED( 173, 11), 
		TO_UNSIGNED( 221, 11), TO_UNSIGNED( 887, 11), TO_UNSIGNED(1041, 11), TO_UNSIGNED(1191, 11), TO_UNSIGNED(1323, 11), TO_UNSIGNED(1792, 11), TO_UNSIGNED( 175, 11), TO_UNSIGNED( 223, 11), 
		TO_UNSIGNED( 890, 11), TO_UNSIGNED(1047, 11), TO_UNSIGNED(1122, 11), TO_UNSIGNED(1335, 11), TO_UNSIGNED(1798, 11), TO_UNSIGNED( 177, 11), TO_UNSIGNED( 225, 11), TO_UNSIGNED( 893, 11), 
		TO_UNSIGNED(1053, 11), TO_UNSIGNED(1125, 11), TO_UNSIGNED(1329, 11), TO_UNSIGNED(1810, 11), TO_UNSIGNED( 179, 11), TO_UNSIGNED( 227, 11), TO_UNSIGNED( 896, 11), TO_UNSIGNED(1059, 11), 
		TO_UNSIGNED(1128, 11), TO_UNSIGNED(1353, 11), TO_UNSIGNED(1786, 11), TO_UNSIGNED(   9, 11), TO_UNSIGNED( 181, 11), TO_UNSIGNED( 229, 11), TO_UNSIGNED( 899, 11), TO_UNSIGNED(1065, 11), 
		TO_UNSIGNED(1131, 11), TO_UNSIGNED(1359, 11), TO_UNSIGNED( 183, 11), TO_UNSIGNED( 231, 11), TO_UNSIGNED( 902, 11), TO_UNSIGNED(1071, 11), TO_UNSIGNED(1134, 11), TO_UNSIGNED(1341, 11), 
		TO_UNSIGNED(1816, 11), TO_UNSIGNED( 139, 11), TO_UNSIGNED( 185, 11), TO_UNSIGNED( 233, 11), TO_UNSIGNED( 905, 11), TO_UNSIGNED(1077, 11), TO_UNSIGNED(1137, 11), TO_UNSIGNED(1347, 11), 
		TO_UNSIGNED( 283, 11), TO_UNSIGNED( 331, 11), TO_UNSIGNED(1000, 11), TO_UNSIGNED(1123, 11), TO_UNSIGNED(1300, 11), TO_UNSIGNED(1616, 11), TO_UNSIGNED(1721, 11), TO_UNSIGNED( 285, 11), 
		TO_UNSIGNED( 333, 11), TO_UNSIGNED(1006, 11), TO_UNSIGNED(1126, 11), TO_UNSIGNED(1294, 11), TO_UNSIGNED(1733, 11), TO_UNSIGNED(1821, 11), TO_UNSIGNED(  14, 11), TO_UNSIGNED( 287, 11), 
		TO_UNSIGNED( 335, 11), TO_UNSIGNED(1012, 11), TO_UNSIGNED(1129, 11), TO_UNSIGNED(1312, 11), TO_UNSIGNED(1727, 11), TO_UNSIGNED(  17, 11), TO_UNSIGNED( 289, 11), TO_UNSIGNED( 337, 11), 
		TO_UNSIGNED(1018, 11), TO_UNSIGNED(1132, 11), TO_UNSIGNED(1306, 11), TO_UNSIGNED(1739, 11), TO_UNSIGNED(  20, 11), TO_UNSIGNED( 291, 11), TO_UNSIGNED( 339, 11), TO_UNSIGNED(1024, 11), 
		TO_UNSIGNED(1135, 11), TO_UNSIGNED(1318, 11), TO_UNSIGNED(1775, 11), TO_UNSIGNED(  23, 11), TO_UNSIGNED( 293, 11), TO_UNSIGNED( 341, 11), TO_UNSIGNED(1030, 11), TO_UNSIGNED(1138, 11), 
		TO_UNSIGNED(1324, 11), TO_UNSIGNED(1781, 11), TO_UNSIGNED(  26, 11), TO_UNSIGNED( 295, 11), TO_UNSIGNED( 343, 11), TO_UNSIGNED(1036, 11), TO_UNSIGNED(1141, 11), TO_UNSIGNED(1336, 11), 
		TO_UNSIGNED(1745, 11), TO_UNSIGNED(  29, 11), TO_UNSIGNED( 297, 11), TO_UNSIGNED( 345, 11), TO_UNSIGNED(1042, 11), TO_UNSIGNED(1144, 11), TO_UNSIGNED(1330, 11), TO_UNSIGNED(1751, 11), 
		TO_UNSIGNED(  32, 11), TO_UNSIGNED( 299, 11), TO_UNSIGNED( 347, 11), TO_UNSIGNED(1048, 11), TO_UNSIGNED(1147, 11), TO_UNSIGNED(1354, 11), TO_UNSIGNED(1757, 11), TO_UNSIGNED(  35, 11), 
		TO_UNSIGNED( 301, 11), TO_UNSIGNED( 349, 11), TO_UNSIGNED(1054, 11), TO_UNSIGNED(1150, 11), TO_UNSIGNED(1360, 11), TO_UNSIGNED(1763, 11), TO_UNSIGNED(  38, 11), TO_UNSIGNED( 303, 11), 
		TO_UNSIGNED( 351, 11), TO_UNSIGNED(1060, 11), TO_UNSIGNED(1153, 11), TO_UNSIGNED(1342, 11), TO_UNSIGNED(1769, 11), TO_UNSIGNED(  41, 11), TO_UNSIGNED( 305, 11), TO_UNSIGNED( 353, 11), 
		TO_UNSIGNED(1066, 11), TO_UNSIGNED(1156, 11), TO_UNSIGNED(1348, 11), TO_UNSIGNED(1805, 11), TO_UNSIGNED(  44, 11), TO_UNSIGNED( 307, 11), TO_UNSIGNED( 355, 11), TO_UNSIGNED(1072, 11), 
		TO_UNSIGNED(1159, 11), TO_UNSIGNED(1372, 11), TO_UNSIGNED(1793, 11), TO_UNSIGNED(  47, 11), TO_UNSIGNED( 309, 11), TO_UNSIGNED( 357, 11), TO_UNSIGNED(1078, 11), TO_UNSIGNED(1162, 11), 
		TO_UNSIGNED(1378, 11), TO_UNSIGNED(1799, 11), TO_UNSIGNED(  50, 11), TO_UNSIGNED( 311, 11), TO_UNSIGNED( 359, 11), TO_UNSIGNED(1084, 11), TO_UNSIGNED(1165, 11), TO_UNSIGNED(1366, 11), 
		TO_UNSIGNED(1811, 11), TO_UNSIGNED(  53, 11), TO_UNSIGNED( 313, 11), TO_UNSIGNED( 361, 11), TO_UNSIGNED(1090, 11), TO_UNSIGNED(1168, 11), TO_UNSIGNED(1396, 11), TO_UNSIGNED(1787, 11), 
		TO_UNSIGNED(  10, 11), TO_UNSIGNED(  56, 11), TO_UNSIGNED( 315, 11), TO_UNSIGNED( 363, 11), TO_UNSIGNED(1096, 11), TO_UNSIGNED(1171, 11), TO_UNSIGNED(1384, 11), TO_UNSIGNED(  59, 11), 
		TO_UNSIGNED( 317, 11), TO_UNSIGNED( 365, 11), TO_UNSIGNED(1102, 11), TO_UNSIGNED(1174, 11), TO_UNSIGNED(1390, 11), TO_UNSIGNED(1817, 11), TO_UNSIGNED(  62, 11), TO_UNSIGNED( 134, 11), 
		TO_UNSIGNED( 140, 11), TO_UNSIGNED( 319, 11), TO_UNSIGNED( 367, 11), TO_UNSIGNED(1108, 11), TO_UNSIGNED(1177, 11), TO_UNSIGNED(  65, 11), TO_UNSIGNED(  82, 11), TO_UNSIGNED( 321, 11), 
		TO_UNSIGNED( 369, 11), TO_UNSIGNED(1114, 11), TO_UNSIGNED(1180, 11), TO_UNSIGNED(1691, 11), TO_UNSIGNED(  68, 11), TO_UNSIGNED( 323, 11), TO_UNSIGNED( 371, 11), TO_UNSIGNED(1120, 11), 
		TO_UNSIGNED(1183, 11), TO_UNSIGNED(1276, 11), TO_UNSIGNED(1715, 11), TO_UNSIGNED(  71, 11), TO_UNSIGNED( 325, 11), TO_UNSIGNED( 373, 11), TO_UNSIGNED( 982, 11), TO_UNSIGNED(1186, 11), 
		TO_UNSIGNED(1282, 11), TO_UNSIGNED(1703, 11), TO_UNSIGNED(  74, 11), TO_UNSIGNED( 327, 11), TO_UNSIGNED( 375, 11), TO_UNSIGNED( 988, 11), TO_UNSIGNED(1189, 11), TO_UNSIGNED(1288, 11), 
		TO_UNSIGNED(1709, 11), TO_UNSIGNED(  77, 11), TO_UNSIGNED( 329, 11), TO_UNSIGNED( 377, 11), TO_UNSIGNED( 994, 11), TO_UNSIGNED(1192, 11), TO_UNSIGNED(1270, 11), TO_UNSIGNED(1697, 11), 
		TO_UNSIGNED( 427, 11), TO_UNSIGNED( 475, 11), TO_UNSIGNED( 944, 11), TO_UNSIGNED(1025, 11), TO_UNSIGNED(1169, 11), TO_UNSIGNED(1343, 11), TO_UNSIGNED(1752, 11), TO_UNSIGNED( 429, 11), 
		TO_UNSIGNED( 477, 11), TO_UNSIGNED( 947, 11), TO_UNSIGNED(1031, 11), TO_UNSIGNED(1172, 11), TO_UNSIGNED(1349, 11), TO_UNSIGNED(1758, 11), TO_UNSIGNED( 431, 11), TO_UNSIGNED( 479, 11), 
		TO_UNSIGNED( 950, 11), TO_UNSIGNED(1037, 11), TO_UNSIGNED(1175, 11), TO_UNSIGNED(1373, 11), TO_UNSIGNED(1764, 11), TO_UNSIGNED( 433, 11), TO_UNSIGNED( 481, 11), TO_UNSIGNED( 953, 11), 
		TO_UNSIGNED(1043, 11), TO_UNSIGNED(1178, 11), TO_UNSIGNED(1379, 11), TO_UNSIGNED(1770, 11), TO_UNSIGNED( 435, 11), TO_UNSIGNED( 483, 11), TO_UNSIGNED( 956, 11), TO_UNSIGNED(1049, 11), 
		TO_UNSIGNED(1181, 11), TO_UNSIGNED(1367, 11), TO_UNSIGNED(1806, 11), TO_UNSIGNED( 437, 11), TO_UNSIGNED( 485, 11), TO_UNSIGNED( 959, 11), TO_UNSIGNED(1055, 11), TO_UNSIGNED(1184, 11), 
		TO_UNSIGNED(1397, 11), TO_UNSIGNED(1794, 11), TO_UNSIGNED( 439, 11), TO_UNSIGNED( 487, 11), TO_UNSIGNED( 962, 11), TO_UNSIGNED(1061, 11), TO_UNSIGNED(1187, 11), TO_UNSIGNED(1385, 11), 
		TO_UNSIGNED(1800, 11), TO_UNSIGNED( 441, 11), TO_UNSIGNED( 489, 11), TO_UNSIGNED( 965, 11), TO_UNSIGNED(1067, 11), TO_UNSIGNED(1190, 11), TO_UNSIGNED(1391, 11), TO_UNSIGNED(1812, 11), 
		TO_UNSIGNED( 135, 11), TO_UNSIGNED( 443, 11), TO_UNSIGNED( 491, 11), TO_UNSIGNED( 968, 11), TO_UNSIGNED(1073, 11), TO_UNSIGNED(1193, 11), TO_UNSIGNED(1788, 11), TO_UNSIGNED(  11, 11), 
		TO_UNSIGNED(  83, 11), TO_UNSIGNED( 445, 11), TO_UNSIGNED( 493, 11), TO_UNSIGNED( 971, 11), TO_UNSIGNED(1079, 11), TO_UNSIGNED(1124, 11), TO_UNSIGNED( 447, 11), TO_UNSIGNED( 495, 11), 
		TO_UNSIGNED( 974, 11), TO_UNSIGNED(1085, 11), TO_UNSIGNED(1127, 11), TO_UNSIGNED(1277, 11), TO_UNSIGNED(1818, 11), TO_UNSIGNED( 141, 11), TO_UNSIGNED( 449, 11), TO_UNSIGNED( 497, 11), 
		TO_UNSIGNED( 977, 11), TO_UNSIGNED(1091, 11), TO_UNSIGNED(1130, 11), TO_UNSIGNED(1283, 11), TO_UNSIGNED( 451, 11), TO_UNSIGNED( 499, 11), TO_UNSIGNED( 908, 11), TO_UNSIGNED(1097, 11), 
		TO_UNSIGNED(1133, 11), TO_UNSIGNED(1289, 11), TO_UNSIGNED(1692, 11), TO_UNSIGNED( 453, 11), TO_UNSIGNED( 501, 11), TO_UNSIGNED( 911, 11), TO_UNSIGNED(1103, 11), TO_UNSIGNED(1136, 11), 
		TO_UNSIGNED(1271, 11), TO_UNSIGNED(1716, 11), TO_UNSIGNED( 455, 11), TO_UNSIGNED( 503, 11), TO_UNSIGNED( 914, 11), TO_UNSIGNED(1109, 11), TO_UNSIGNED(1139, 11), TO_UNSIGNED(1301, 11), 
		TO_UNSIGNED(1704, 11), TO_UNSIGNED( 457, 11), TO_UNSIGNED( 505, 11), TO_UNSIGNED( 917, 11), TO_UNSIGNED(1115, 11), TO_UNSIGNED(1142, 11), TO_UNSIGNED(1295, 11), TO_UNSIGNED(1710, 11), 
		TO_UNSIGNED( 459, 11), TO_UNSIGNED( 507, 11), TO_UNSIGNED( 920, 11), TO_UNSIGNED(1121, 11), TO_UNSIGNED(1145, 11), TO_UNSIGNED(1313, 11), TO_UNSIGNED(1698, 11), TO_UNSIGNED( 461, 11), 
		TO_UNSIGNED( 509, 11), TO_UNSIGNED( 923, 11), TO_UNSIGNED( 983, 11), TO_UNSIGNED(1148, 11), TO_UNSIGNED(1307, 11), TO_UNSIGNED(1722, 11), TO_UNSIGNED( 463, 11), TO_UNSIGNED( 511, 11), 
		TO_UNSIGNED( 926, 11), TO_UNSIGNED( 989, 11), TO_UNSIGNED(1151, 11), TO_UNSIGNED(1319, 11), TO_UNSIGNED(1734, 11), TO_UNSIGNED( 465, 11), TO_UNSIGNED( 513, 11), TO_UNSIGNED( 929, 11), 
		TO_UNSIGNED( 995, 11), TO_UNSIGNED(1154, 11), TO_UNSIGNED(1325, 11), TO_UNSIGNED(1728, 11), TO_UNSIGNED( 467, 11), TO_UNSIGNED( 515, 11), TO_UNSIGNED( 932, 11), TO_UNSIGNED(1001, 11), 
		TO_UNSIGNED(1157, 11), TO_UNSIGNED(1337, 11), TO_UNSIGNED(1740, 11), TO_UNSIGNED( 469, 11), TO_UNSIGNED( 517, 11), TO_UNSIGNED( 935, 11), TO_UNSIGNED(1007, 11), TO_UNSIGNED(1160, 11), 
		TO_UNSIGNED(1331, 11), TO_UNSIGNED(1776, 11), TO_UNSIGNED( 471, 11), TO_UNSIGNED( 519, 11), TO_UNSIGNED( 938, 11), TO_UNSIGNED(1013, 11), TO_UNSIGNED(1163, 11), TO_UNSIGNED(1355, 11), 
		TO_UNSIGNED(1782, 11), TO_UNSIGNED( 473, 11), TO_UNSIGNED( 521, 11), TO_UNSIGNED( 941, 11), TO_UNSIGNED(1019, 11), TO_UNSIGNED(1166, 11), TO_UNSIGNED(1361, 11), TO_UNSIGNED(1746, 11)
	);                        

	SIGNAL  READ_C : UNSIGNED(10 downto 0);
	SIGNAL WRITE_C : UNSIGNED(10 downto 0);
	SIGNAL ROM_ADR : UNSIGNED(10 downto 0);

	SIGNAL IN_BIS : STD_LOGIC_VECTOR (15 downto 0);
	SIGNAL WE_BIS : STD_LOGIC;
	
BEGIN

	-------------------------------------------------------------------------
	-- synthesis translate_off 
  	PROCESS
  	BEGIN
    	WAIT FOR 1 ns;
		printmsg("(IMS) Q16_8_C_to_V_RAM : ALLOCATION OK !");
    	WAIT;
  	END PROCESS;
	-- synthesis translate_on 
	-------------------------------------------------------------------------

	--
	--
	--
	PROCESS(clock, reset)
		VARIABLE TEMP : UNSIGNED(10 downto 0);
	BEGIN
		IF reset = '0' THEN
			WRITE_C <= TO_UNSIGNED(0, 11);
		elsif clock'event and clock = '1' THEN
			IF WRITE_EN = '1' AND HOLDN = '1' THEN
				TEMP := WRITE_C + TO_UNSIGNED(1, 11);
				IF TEMP = 1824 THEN
					TEMP := TO_UNSIGNED(0, 11);
				END IF;
				WE_BIS  <= '1';
				WRITE_C <= TEMP;
			ELSE
				WE_BIS  <= '0';
				WRITE_C <= WRITE_C;
			END IF;
			IN_BIS  <= INPUT_1(15 downto 0);
		END if;
	END PROCESS;


	--
	--
	--
	process(clock, reset)
		VARIABLE TEMP : UNSIGNED(10 downto 0);
		VARIABLE TMP  : STD_LOGIC_VECTOR(15 downto 0);
	begin
		if reset = '0' then
			READ_C  <= TO_UNSIGNED(0, 11);
		elsif clock'event and clock = '1' then
			TEMP := READ_C;
			if read_en = '1' AND holdn = '1' then
				TEMP := TEMP + TO_UNSIGNED(1, 11);
				IF TEMP = 1824 THEN
					TEMP := TO_UNSIGNED(0, 11);
				END IF;
			end if;
			READ_C <= TEMP;
			TMP := RAM( to_integer( TEMP ) );
			OUTPUT_1 <= STD_LOGIC_VECTOR(RESIZE( SIGNED( TMP ), 32 )) ;
		end if;
	end process;


	--
	--
	--
	process(clock)
		VARIABLE ADR : INTEGER RANGE 0 to 1823;
		VARIABLE POS : INTEGER RANGE 0 to 1823;
	begin
		if clock'event and clock = '1' then
			ADR     := to_integer( WRITE_C );
			ROM_ADR <= ROM( ADR );
		end if;
	end process;


	--
	--
	--
	process(clock)
		VARIABLE TMP : STD_LOGIC_VECTOR(15 downto 0);
	begin
--		IF reset = '0' THEN
--				OUTPUT_1 <= (OTHERS => '0');
		if clock'event and clock = '1' then
			if WE_BIS = '1' then
	-- synthesis translate_off 
	--			printmsg("(Q16_8_V_to_C_RAM) ===> WRITING (" & to_int_str( STD_LOGIC_VECTOR(IN_BIS),6) & ") AT POSITION : " & to_int_str( STD_LOGIC_VECTOR(ROM_ADR),6) );
	-- synthesis translate_on
				RAM( to_integer( ROM_ADR ) ) <= IN_BIS;
			end if;
		end if;
	end process;
	
END cRAM;
