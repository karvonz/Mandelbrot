library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------
-- synthesis translate_off 
--library ims;
--use ims.coprocessor.all;
-- synthesis translate_on 
-------------------------------------------------------------------------

ENTITY Q16_8_IndexRAM is
	PORT (
		RESET    : in  STD_LOGIC;
		CLOCK    : in  STD_LOGIC;
		WRITE_EN : in  STD_LOGIC;
		READ_EN  : in  STD_LOGIC;
		INPUT_1  : in  STD_LOGIC_VECTOR(15 downto 0);
		OUTPUT_1 : out STD_LOGIC_VECTOR(15 downto 0)
	);
END;

architecture cRAM of Q16_8_IndexRAM is
   type ram_type is array (0 to 1824-1) of STD_LOGIC_VECTOR (15 downto 0);                 
   type rom_type is array (0 to 1824-1) of UNSIGNED (11 downto 0);                 
   signal RAM : ram_type;

   signal WE_BIS : STD_LOGIC;
   signal IN_BIS : STD_LOGIC_VECTOR (15 downto 0);

   constant ROM : rom_type:= (
		TO_UNSIGNED(75, 12),   TO_UNSIGNED(618, 12), 
		TO_UNSIGNED(732, 12),  TO_UNSIGNED(1425, 12), 
		TO_UNSIGNED(1500, 12), TO_UNSIGNED(1683, 12), 
		TO_UNSIGNED(84, 12),   TO_UNSIGNED(621, 12), 
		TO_UNSIGNED(738, 12),  TO_UNSIGNED(1428, 12), 
		TO_UNSIGNED(1506, 12), TO_UNSIGNED(1614, 12), 
		TO_UNSIGNED(86, 12),   TO_UNSIGNED(624, 12), 
		TO_UNSIGNED(744, 12),  TO_UNSIGNED(1437, 12), 
		TO_UNSIGNED(1488, 12), TO_UNSIGNED(1819, 12), 
		TO_UNSIGNED(12, 12),   TO_UNSIGNED(88, 12), 
		TO_UNSIGNED(627, 12),  TO_UNSIGNED(750, 12), 
		TO_UNSIGNED(1440, 12), TO_UNSIGNED(1512, 12), 
		TO_UNSIGNED(15, 12),   TO_UNSIGNED(90, 12), 
		TO_UNSIGNED(630, 12),  TO_UNSIGNED(756, 12), 
		TO_UNSIGNED(1443, 12), TO_UNSIGNED(1524, 12), 
		TO_UNSIGNED(18, 12),   TO_UNSIGNED(92, 12), 
		TO_UNSIGNED(633, 12),  TO_UNSIGNED(762, 12), 
		TO_UNSIGNED(1446, 12), TO_UNSIGNED(1518, 12), 
		TO_UNSIGNED(21, 12),   TO_UNSIGNED(94, 12), 
		TO_UNSIGNED(636, 12), TO_UNSIGNED(768, 12), 
  TO_UNSIGNED(1449, 12), TO_UNSIGNED(1542, 12), 
  TO_UNSIGNED(24, 12), TO_UNSIGNED(96, 12), 
  TO_UNSIGNED(639, 12), TO_UNSIGNED(774, 12), 
  TO_UNSIGNED(1452, 12), TO_UNSIGNED(1548, 12), 
  TO_UNSIGNED(27, 12), TO_UNSIGNED(98, 12), 
  TO_UNSIGNED(642, 12), TO_UNSIGNED(780, 12), 
  TO_UNSIGNED(1455, 12), TO_UNSIGNED(1530, 12), 
  TO_UNSIGNED(30, 12), TO_UNSIGNED(100, 12), 
  TO_UNSIGNED(645, 12), TO_UNSIGNED(786, 12), 
  TO_UNSIGNED(1461, 12), TO_UNSIGNED(1536, 12), 
  TO_UNSIGNED(33, 12), TO_UNSIGNED(102, 12), 
  TO_UNSIGNED(648, 12), TO_UNSIGNED(792, 12), 
  TO_UNSIGNED(1458, 12), TO_UNSIGNED(1554, 12), 
  TO_UNSIGNED(36, 12), TO_UNSIGNED(104, 12), 
  TO_UNSIGNED(651, 12), TO_UNSIGNED(798, 12), 
  TO_UNSIGNED(1485, 12), TO_UNSIGNED(1560, 12), 
  TO_UNSIGNED(39, 12), TO_UNSIGNED(106, 12), 
  TO_UNSIGNED(654, 12), TO_UNSIGNED(804, 12), 
  TO_UNSIGNED(1572, 12), TO_UNSIGNED(1617, 12), 
  TO_UNSIGNED(42, 12), TO_UNSIGNED(108, 12), 
  TO_UNSIGNED(657, 12), TO_UNSIGNED(810, 12), 
  TO_UNSIGNED(1398, 12), TO_UNSIGNED(1566, 12), 
  TO_UNSIGNED(45, 12), TO_UNSIGNED(110, 12), 
  TO_UNSIGNED(660, 12), TO_UNSIGNED(816, 12), 
  TO_UNSIGNED(1401, 12), TO_UNSIGNED(1584, 12), 
  TO_UNSIGNED(48, 12), TO_UNSIGNED(112, 12), 
  TO_UNSIGNED(663, 12), TO_UNSIGNED(822, 12), 
  TO_UNSIGNED(1404, 12), TO_UNSIGNED(1578, 12), 
  TO_UNSIGNED(51, 12), TO_UNSIGNED(114, 12), 
  TO_UNSIGNED(666, 12), TO_UNSIGNED(828, 12), 
  TO_UNSIGNED(1413, 12), TO_UNSIGNED(1596, 12), 
  TO_UNSIGNED(54, 12), TO_UNSIGNED(116, 12), 
  TO_UNSIGNED(669, 12), TO_UNSIGNED(690, 12), 
  TO_UNSIGNED(1416, 12), TO_UNSIGNED(1602, 12), 
  TO_UNSIGNED(57, 12), TO_UNSIGNED(118, 12), 
  TO_UNSIGNED(672, 12), TO_UNSIGNED(696, 12), 
  TO_UNSIGNED(1419, 12), TO_UNSIGNED(1590, 12), 
  TO_UNSIGNED(0, 12), TO_UNSIGNED(60, 12), 
  TO_UNSIGNED(120, 12), TO_UNSIGNED(675, 12), 
  TO_UNSIGNED(702, 12), TO_UNSIGNED(1407, 12), 
  TO_UNSIGNED(63, 12), TO_UNSIGNED(122, 12), 
  TO_UNSIGNED(678, 12), TO_UNSIGNED(708, 12), 
  TO_UNSIGNED(1410, 12), TO_UNSIGNED(1476, 12), 
  TO_UNSIGNED(66, 12), TO_UNSIGNED(124, 12), 
  TO_UNSIGNED(681, 12), TO_UNSIGNED(714, 12), 
  TO_UNSIGNED(1434, 12), TO_UNSIGNED(1464, 12), 
  TO_UNSIGNED(69, 12), TO_UNSIGNED(126, 12), 
  TO_UNSIGNED(684, 12), TO_UNSIGNED(720, 12), 
  TO_UNSIGNED(1431, 12), TO_UNSIGNED(1470, 12), 
  TO_UNSIGNED(72, 12), TO_UNSIGNED(128, 12), 
  TO_UNSIGNED(687, 12), TO_UNSIGNED(726, 12), 
  TO_UNSIGNED(1422, 12), TO_UNSIGNED(1494, 12), 
  TO_UNSIGNED(186, 12), TO_UNSIGNED(234, 12), 
  TO_UNSIGNED(775, 12), TO_UNSIGNED(906, 12), 
  TO_UNSIGNED(1435, 12), TO_UNSIGNED(1585, 12), 
  TO_UNSIGNED(188, 12), TO_UNSIGNED(236, 12), 
  TO_UNSIGNED(781, 12), TO_UNSIGNED(909, 12), 
  TO_UNSIGNED(1432, 12), TO_UNSIGNED(1579, 12), 
  TO_UNSIGNED(190, 12), TO_UNSIGNED(238, 12), 
  TO_UNSIGNED(787, 12), TO_UNSIGNED(912, 12), 
  TO_UNSIGNED(1423, 12), TO_UNSIGNED(1597, 12), 
  TO_UNSIGNED(192, 12), TO_UNSIGNED(240, 12), 
  TO_UNSIGNED(793, 12), TO_UNSIGNED(915, 12), 
  TO_UNSIGNED(1426, 12), TO_UNSIGNED(1603, 12), 
  TO_UNSIGNED(194, 12), TO_UNSIGNED(242, 12), 
  TO_UNSIGNED(799, 12), TO_UNSIGNED(918, 12), 
  TO_UNSIGNED(1429, 12), TO_UNSIGNED(1591, 12), 
  TO_UNSIGNED(1, 12), TO_UNSIGNED(196, 12), 
  TO_UNSIGNED(244, 12), TO_UNSIGNED(805, 12), 
  TO_UNSIGNED(921, 12), TO_UNSIGNED(1438, 12), 
  TO_UNSIGNED(198, 12), TO_UNSIGNED(246, 12), 
  TO_UNSIGNED(811, 12), TO_UNSIGNED(924, 12), 
  TO_UNSIGNED(1441, 12), TO_UNSIGNED(1477, 12), 
  TO_UNSIGNED(200, 12), TO_UNSIGNED(248, 12), 
  TO_UNSIGNED(817, 12), TO_UNSIGNED(927, 12), 
  TO_UNSIGNED(1444, 12), TO_UNSIGNED(1465, 12), 
  TO_UNSIGNED(202, 12), TO_UNSIGNED(250, 12), 
  TO_UNSIGNED(823, 12), TO_UNSIGNED(930, 12), 
  TO_UNSIGNED(1447, 12), TO_UNSIGNED(1471, 12), 
  TO_UNSIGNED(204, 12), TO_UNSIGNED(252, 12), 
  TO_UNSIGNED(829, 12), TO_UNSIGNED(933, 12), 
  TO_UNSIGNED(1450, 12), TO_UNSIGNED(1495, 12), 
  TO_UNSIGNED(206, 12), TO_UNSIGNED(254, 12), 
  TO_UNSIGNED(691, 12), TO_UNSIGNED(936, 12), 
  TO_UNSIGNED(1453, 12), TO_UNSIGNED(1501, 12), 
  TO_UNSIGNED(208, 12), TO_UNSIGNED(256, 12), 
  TO_UNSIGNED(697, 12), TO_UNSIGNED(939, 12), 
  TO_UNSIGNED(1456, 12), TO_UNSIGNED(1507, 12), 
  TO_UNSIGNED(210, 12), TO_UNSIGNED(258, 12), 
  TO_UNSIGNED(703, 12), TO_UNSIGNED(942, 12), 
  TO_UNSIGNED(1462, 12), TO_UNSIGNED(1489, 12), 
  TO_UNSIGNED(212, 12), TO_UNSIGNED(260, 12), 
  TO_UNSIGNED(709, 12), TO_UNSIGNED(945, 12), 
  TO_UNSIGNED(1459, 12), TO_UNSIGNED(1513, 12), 
  TO_UNSIGNED(214, 12), TO_UNSIGNED(262, 12), 
  TO_UNSIGNED(715, 12), TO_UNSIGNED(948, 12), 
  TO_UNSIGNED(1486, 12), TO_UNSIGNED(1525, 12), 
  TO_UNSIGNED(216, 12), TO_UNSIGNED(264, 12), 
  TO_UNSIGNED(721, 12), TO_UNSIGNED(951, 12), 
  TO_UNSIGNED(1519, 12), TO_UNSIGNED(1618, 12), 
  TO_UNSIGNED(218, 12), TO_UNSIGNED(266, 12), 
  TO_UNSIGNED(727, 12), TO_UNSIGNED(954, 12), 
  TO_UNSIGNED(1399, 12), TO_UNSIGNED(1543, 12), 
  TO_UNSIGNED(220, 12), TO_UNSIGNED(268, 12), 
  TO_UNSIGNED(733, 12), TO_UNSIGNED(957, 12), 
  TO_UNSIGNED(1402, 12), TO_UNSIGNED(1549, 12), 
  TO_UNSIGNED(222, 12), TO_UNSIGNED(270, 12), 
  TO_UNSIGNED(739, 12), TO_UNSIGNED(960, 12), 
  TO_UNSIGNED(1405, 12), TO_UNSIGNED(1531, 12), 
  TO_UNSIGNED(224, 12), TO_UNSIGNED(272, 12), 
  TO_UNSIGNED(745, 12), TO_UNSIGNED(963, 12), 
  TO_UNSIGNED(1414, 12), TO_UNSIGNED(1537, 12), 
  TO_UNSIGNED(226, 12), TO_UNSIGNED(274, 12), 
  TO_UNSIGNED(751, 12), TO_UNSIGNED(966, 12), 
  TO_UNSIGNED(1417, 12), TO_UNSIGNED(1555, 12), 
  TO_UNSIGNED(228, 12), TO_UNSIGNED(276, 12), 
  TO_UNSIGNED(757, 12), TO_UNSIGNED(969, 12), 
  TO_UNSIGNED(1420, 12), TO_UNSIGNED(1561, 12), 
  TO_UNSIGNED(230, 12), TO_UNSIGNED(278, 12), 
  TO_UNSIGNED(763, 12), TO_UNSIGNED(972, 12), 
  TO_UNSIGNED(1408, 12), TO_UNSIGNED(1573, 12), 
  TO_UNSIGNED(232, 12), TO_UNSIGNED(280, 12), 
  TO_UNSIGNED(769, 12), TO_UNSIGNED(975, 12), 
  TO_UNSIGNED(1411, 12), TO_UNSIGNED(1567, 12), 
  TO_UNSIGNED(235, 12), TO_UNSIGNED(282, 12), 
  TO_UNSIGNED(788, 12), TO_UNSIGNED(1206, 12), 
  TO_UNSIGNED(1556, 12), TO_UNSIGNED(1635, 12), 
  TO_UNSIGNED(237, 12), TO_UNSIGNED(284, 12), 
  TO_UNSIGNED(794, 12), TO_UNSIGNED(1209, 12), 
  TO_UNSIGNED(1562, 12), TO_UNSIGNED(1629, 12), 
  TO_UNSIGNED(239, 12), TO_UNSIGNED(286, 12), 
  TO_UNSIGNED(800, 12), TO_UNSIGNED(1194, 12), 
  TO_UNSIGNED(1574, 12), TO_UNSIGNED(1632, 12), 
  TO_UNSIGNED(241, 12), TO_UNSIGNED(288, 12), 
  TO_UNSIGNED(806, 12), TO_UNSIGNED(1215, 12), 
  TO_UNSIGNED(1568, 12), TO_UNSIGNED(1641, 12), 
  TO_UNSIGNED(243, 12), TO_UNSIGNED(290, 12), 
  TO_UNSIGNED(812, 12), TO_UNSIGNED(1212, 12), 
  TO_UNSIGNED(1586, 12), TO_UNSIGNED(1638, 12), 
  TO_UNSIGNED(245, 12), TO_UNSIGNED(292, 12), 
  TO_UNSIGNED(818, 12), TO_UNSIGNED(1221, 12), 
  TO_UNSIGNED(1580, 12), TO_UNSIGNED(1644, 12), 
  TO_UNSIGNED(247, 12), TO_UNSIGNED(294, 12), 
  TO_UNSIGNED(824, 12), TO_UNSIGNED(1224, 12), 
  TO_UNSIGNED(1598, 12), TO_UNSIGNED(1650, 12), 
  TO_UNSIGNED(249, 12), TO_UNSIGNED(296, 12), 
  TO_UNSIGNED(830, 12), TO_UNSIGNED(1227, 12), 
  TO_UNSIGNED(1604, 12), TO_UNSIGNED(1647, 12), 
  TO_UNSIGNED(251, 12), TO_UNSIGNED(298, 12), 
  TO_UNSIGNED(692, 12), TO_UNSIGNED(1218, 12), 
  TO_UNSIGNED(1592, 12), TO_UNSIGNED(1653, 12), 
  TO_UNSIGNED(2, 12), TO_UNSIGNED(253, 12), 
  TO_UNSIGNED(300, 12), TO_UNSIGNED(698, 12), 
  TO_UNSIGNED(1233, 12), TO_UNSIGNED(1656, 12), 
  TO_UNSIGNED(255, 12), TO_UNSIGNED(302, 12), 
  TO_UNSIGNED(704, 12), TO_UNSIGNED(1236, 12), 
  TO_UNSIGNED(1478, 12), TO_UNSIGNED(1659, 12), 
  TO_UNSIGNED(257, 12), TO_UNSIGNED(304, 12), 
  TO_UNSIGNED(710, 12), TO_UNSIGNED(1239, 12), 
  TO_UNSIGNED(1466, 12), TO_UNSIGNED(1662, 12), 
  TO_UNSIGNED(259, 12), TO_UNSIGNED(306, 12), 
  TO_UNSIGNED(716, 12), TO_UNSIGNED(1230, 12), 
  TO_UNSIGNED(1472, 12), TO_UNSIGNED(1665, 12), 
  TO_UNSIGNED(261, 12), TO_UNSIGNED(308, 12), 
  TO_UNSIGNED(722, 12), TO_UNSIGNED(1251, 12), 
  TO_UNSIGNED(1496, 12), TO_UNSIGNED(1671, 12), 
  TO_UNSIGNED(263, 12), TO_UNSIGNED(310, 12), 
  TO_UNSIGNED(728, 12), TO_UNSIGNED(1242, 12), 
  TO_UNSIGNED(1502, 12), TO_UNSIGNED(1668, 12), 
  TO_UNSIGNED(265, 12), TO_UNSIGNED(312, 12), 
  TO_UNSIGNED(734, 12), TO_UNSIGNED(1245, 12), 
  TO_UNSIGNED(1508, 12), TO_UNSIGNED(1674, 12), 
  TO_UNSIGNED(267, 12), TO_UNSIGNED(314, 12), 
  TO_UNSIGNED(740, 12), TO_UNSIGNED(1248, 12), 
  TO_UNSIGNED(1490, 12), TO_UNSIGNED(1677, 12), 
  TO_UNSIGNED(269, 12), TO_UNSIGNED(316, 12), 
  TO_UNSIGNED(746, 12), TO_UNSIGNED(1257, 12), 
  TO_UNSIGNED(1514, 12), TO_UNSIGNED(1680, 12), 
  TO_UNSIGNED(271, 12), TO_UNSIGNED(318, 12), 
  TO_UNSIGNED(752, 12), TO_UNSIGNED(1254, 12), 
  TO_UNSIGNED(1482, 12), TO_UNSIGNED(1526, 12), 
  TO_UNSIGNED(273, 12), TO_UNSIGNED(320, 12), 
  TO_UNSIGNED(758, 12), TO_UNSIGNED(1263, 12), 
  TO_UNSIGNED(1520, 12), TO_UNSIGNED(1608, 12), 
  TO_UNSIGNED(275, 12), TO_UNSIGNED(322, 12), 
  TO_UNSIGNED(764, 12), TO_UNSIGNED(1260, 12), 
  TO_UNSIGNED(1544, 12), TO_UNSIGNED(1611, 12), 
  TO_UNSIGNED(277, 12), TO_UNSIGNED(324, 12), 
  TO_UNSIGNED(770, 12), TO_UNSIGNED(1197, 12), 
  TO_UNSIGNED(1550, 12), TO_UNSIGNED(1620, 12), 
  TO_UNSIGNED(279, 12), TO_UNSIGNED(326, 12), 
  TO_UNSIGNED(776, 12), TO_UNSIGNED(1200, 12), 
  TO_UNSIGNED(1532, 12), TO_UNSIGNED(1623, 12), 
  TO_UNSIGNED(281, 12), TO_UNSIGNED(328, 12), 
  TO_UNSIGNED(782, 12), TO_UNSIGNED(1203, 12), 
  TO_UNSIGNED(1538, 12), TO_UNSIGNED(1626, 12), 
  TO_UNSIGNED(330, 12), TO_UNSIGNED(378, 12), 
  TO_UNSIGNED(705, 12), TO_UNSIGNED(885, 12), 
  TO_UNSIGNED(1605, 12), TO_UNSIGNED(1669, 12), 
  TO_UNSIGNED(332, 12), TO_UNSIGNED(380, 12), 
  TO_UNSIGNED(711, 12), TO_UNSIGNED(888, 12), 
  TO_UNSIGNED(1593, 12), TO_UNSIGNED(1675, 12), 
  TO_UNSIGNED(3, 12), TO_UNSIGNED(334, 12), 
  TO_UNSIGNED(382, 12), TO_UNSIGNED(717, 12), 
  TO_UNSIGNED(891, 12), TO_UNSIGNED(1678, 12), 
  TO_UNSIGNED(336, 12), TO_UNSIGNED(384, 12), 
  TO_UNSIGNED(723, 12), TO_UNSIGNED(894, 12), 
  TO_UNSIGNED(1479, 12), TO_UNSIGNED(1681, 12), 
  TO_UNSIGNED(338, 12), TO_UNSIGNED(386, 12), 
  TO_UNSIGNED(729, 12), TO_UNSIGNED(897, 12), 
  TO_UNSIGNED(1467, 12), TO_UNSIGNED(1483, 12), 
  TO_UNSIGNED(340, 12), TO_UNSIGNED(388, 12), 
  TO_UNSIGNED(735, 12), TO_UNSIGNED(900, 12), 
  TO_UNSIGNED(1473, 12), TO_UNSIGNED(1609, 12), 
  TO_UNSIGNED(342, 12), TO_UNSIGNED(390, 12), 
  TO_UNSIGNED(741, 12), TO_UNSIGNED(903, 12), 
  TO_UNSIGNED(1497, 12), TO_UNSIGNED(1612, 12), 
  TO_UNSIGNED(344, 12), TO_UNSIGNED(392, 12), 
  TO_UNSIGNED(747, 12), TO_UNSIGNED(834, 12), 
  TO_UNSIGNED(1503, 12), TO_UNSIGNED(1621, 12), 
  TO_UNSIGNED(346, 12), TO_UNSIGNED(394, 12), 
  TO_UNSIGNED(753, 12), TO_UNSIGNED(837, 12), 
  TO_UNSIGNED(1509, 12), TO_UNSIGNED(1624, 12), 
  TO_UNSIGNED(348, 12), TO_UNSIGNED(396, 12), 
  TO_UNSIGNED(759, 12), TO_UNSIGNED(840, 12), 
  TO_UNSIGNED(1491, 12), TO_UNSIGNED(1627, 12), 
  TO_UNSIGNED(350, 12), TO_UNSIGNED(398, 12), 
  TO_UNSIGNED(765, 12), TO_UNSIGNED(843, 12), 
  TO_UNSIGNED(1515, 12), TO_UNSIGNED(1636, 12), 
  TO_UNSIGNED(352, 12), TO_UNSIGNED(400, 12), 
  TO_UNSIGNED(771, 12), TO_UNSIGNED(846, 12), 
  TO_UNSIGNED(1527, 12), TO_UNSIGNED(1630, 12), 
  TO_UNSIGNED(354, 12), TO_UNSIGNED(402, 12), 
  TO_UNSIGNED(777, 12), TO_UNSIGNED(849, 12), 
  TO_UNSIGNED(1521, 12), TO_UNSIGNED(1633, 12), 
  TO_UNSIGNED(356, 12), TO_UNSIGNED(404, 12), 
  TO_UNSIGNED(783, 12), TO_UNSIGNED(852, 12), 
  TO_UNSIGNED(1545, 12), TO_UNSIGNED(1642, 12), 
  TO_UNSIGNED(358, 12), TO_UNSIGNED(406, 12), 
  TO_UNSIGNED(789, 12), TO_UNSIGNED(855, 12), 
  TO_UNSIGNED(1551, 12), TO_UNSIGNED(1639, 12), 
  TO_UNSIGNED(360, 12), TO_UNSIGNED(408, 12), 
  TO_UNSIGNED(795, 12), TO_UNSIGNED(858, 12), 
  TO_UNSIGNED(1533, 12), TO_UNSIGNED(1645, 12), 
  TO_UNSIGNED(362, 12), TO_UNSIGNED(410, 12), 
  TO_UNSIGNED(801, 12), TO_UNSIGNED(861, 12), 
  TO_UNSIGNED(1539, 12), TO_UNSIGNED(1651, 12), 
  TO_UNSIGNED(364, 12), TO_UNSIGNED(412, 12), 
  TO_UNSIGNED(807, 12), TO_UNSIGNED(864, 12), 
  TO_UNSIGNED(1557, 12), TO_UNSIGNED(1648, 12), 
  TO_UNSIGNED(366, 12), TO_UNSIGNED(414, 12), 
  TO_UNSIGNED(813, 12), TO_UNSIGNED(867, 12), 
  TO_UNSIGNED(1563, 12), TO_UNSIGNED(1654, 12), 
  TO_UNSIGNED(368, 12), TO_UNSIGNED(416, 12), 
  TO_UNSIGNED(819, 12), TO_UNSIGNED(870, 12), 
  TO_UNSIGNED(1575, 12), TO_UNSIGNED(1657, 12), 
  TO_UNSIGNED(370, 12), TO_UNSIGNED(418, 12), 
  TO_UNSIGNED(825, 12), TO_UNSIGNED(873, 12), 
  TO_UNSIGNED(1569, 12), TO_UNSIGNED(1660, 12), 
  TO_UNSIGNED(372, 12), TO_UNSIGNED(420, 12), 
  TO_UNSIGNED(831, 12), TO_UNSIGNED(876, 12), 
  TO_UNSIGNED(1587, 12), TO_UNSIGNED(1663, 12), 
  TO_UNSIGNED(374, 12), TO_UNSIGNED(422, 12), 
  TO_UNSIGNED(693, 12), TO_UNSIGNED(879, 12), 
  TO_UNSIGNED(1581, 12), TO_UNSIGNED(1666, 12), 
  TO_UNSIGNED(376, 12), TO_UNSIGNED(424, 12), 
  TO_UNSIGNED(699, 12), TO_UNSIGNED(882, 12), 
  TO_UNSIGNED(1599, 12), TO_UNSIGNED(1672, 12), 
  TO_UNSIGNED(379, 12), TO_UNSIGNED(426, 12), 
  TO_UNSIGNED(682, 12), TO_UNSIGNED(736, 12), 
  TO_UNSIGNED(1198, 12), TO_UNSIGNED(1540, 12), 
  TO_UNSIGNED(381, 12), TO_UNSIGNED(428, 12), 
  TO_UNSIGNED(685, 12), TO_UNSIGNED(742, 12), 
  TO_UNSIGNED(1201, 12), TO_UNSIGNED(1558, 12), 
  TO_UNSIGNED(383, 12), TO_UNSIGNED(430, 12), 
  TO_UNSIGNED(688, 12), TO_UNSIGNED(748, 12), 
  TO_UNSIGNED(1204, 12), TO_UNSIGNED(1564, 12), 
  TO_UNSIGNED(385, 12), TO_UNSIGNED(432, 12), 
  TO_UNSIGNED(619, 12), TO_UNSIGNED(754, 12), 
  TO_UNSIGNED(1207, 12), TO_UNSIGNED(1576, 12), 
  TO_UNSIGNED(387, 12), TO_UNSIGNED(434, 12), 
  TO_UNSIGNED(622, 12), TO_UNSIGNED(760, 12), 
  TO_UNSIGNED(1210, 12), TO_UNSIGNED(1570, 12), 
  TO_UNSIGNED(389, 12), TO_UNSIGNED(436, 12), 
  TO_UNSIGNED(625, 12), TO_UNSIGNED(766, 12), 
  TO_UNSIGNED(1195, 12), TO_UNSIGNED(1588, 12), 
  TO_UNSIGNED(391, 12), TO_UNSIGNED(438, 12), 
  TO_UNSIGNED(628, 12), TO_UNSIGNED(772, 12), 
  TO_UNSIGNED(1216, 12), TO_UNSIGNED(1582, 12), 
  TO_UNSIGNED(393, 12), TO_UNSIGNED(440, 12), 
  TO_UNSIGNED(631, 12), TO_UNSIGNED(778, 12), 
  TO_UNSIGNED(1213, 12), TO_UNSIGNED(1600, 12), 
  TO_UNSIGNED(395, 12), TO_UNSIGNED(442, 12), 
  TO_UNSIGNED(634, 12), TO_UNSIGNED(784, 12), 
  TO_UNSIGNED(1222, 12), TO_UNSIGNED(1606, 12), 
  TO_UNSIGNED(397, 12), TO_UNSIGNED(444, 12), 
  TO_UNSIGNED(637, 12), TO_UNSIGNED(790, 12), 
  TO_UNSIGNED(1225, 12), TO_UNSIGNED(1594, 12), 
  TO_UNSIGNED(4, 12), TO_UNSIGNED(399, 12), 
  TO_UNSIGNED(446, 12), TO_UNSIGNED(640, 12), 
  TO_UNSIGNED(796, 12), TO_UNSIGNED(1228, 12), 
  TO_UNSIGNED(401, 12), TO_UNSIGNED(448, 12), 
  TO_UNSIGNED(643, 12), TO_UNSIGNED(802, 12), 
  TO_UNSIGNED(1219, 12), TO_UNSIGNED(1480, 12), 
  TO_UNSIGNED(403, 12), TO_UNSIGNED(450, 12), 
  TO_UNSIGNED(646, 12), TO_UNSIGNED(808, 12), 
  TO_UNSIGNED(1234, 12), TO_UNSIGNED(1468, 12), 
  TO_UNSIGNED(405, 12), TO_UNSIGNED(452, 12), 
  TO_UNSIGNED(649, 12), TO_UNSIGNED(814, 12), 
  TO_UNSIGNED(1237, 12), TO_UNSIGNED(1474, 12), 
  TO_UNSIGNED(407, 12), TO_UNSIGNED(454, 12), 
  TO_UNSIGNED(652, 12), TO_UNSIGNED(820, 12), 
  TO_UNSIGNED(1240, 12), TO_UNSIGNED(1498, 12), 
  TO_UNSIGNED(409, 12), TO_UNSIGNED(456, 12), 
  TO_UNSIGNED(655, 12), TO_UNSIGNED(826, 12), 
  TO_UNSIGNED(1231, 12), TO_UNSIGNED(1504, 12), 
  TO_UNSIGNED(411, 12), TO_UNSIGNED(458, 12), 
  TO_UNSIGNED(658, 12), TO_UNSIGNED(832, 12), 
  TO_UNSIGNED(1252, 12), TO_UNSIGNED(1510, 12), 
  TO_UNSIGNED(413, 12), TO_UNSIGNED(460, 12), 
  TO_UNSIGNED(661, 12), TO_UNSIGNED(694, 12), 
  TO_UNSIGNED(1243, 12), TO_UNSIGNED(1492, 12), 
  TO_UNSIGNED(415, 12), TO_UNSIGNED(462, 12), 
  TO_UNSIGNED(664, 12), TO_UNSIGNED(700, 12), 
  TO_UNSIGNED(1246, 12), TO_UNSIGNED(1516, 12), 
  TO_UNSIGNED(417, 12), TO_UNSIGNED(464, 12), 
  TO_UNSIGNED(667, 12), TO_UNSIGNED(706, 12), 
  TO_UNSIGNED(1249, 12), TO_UNSIGNED(1528, 12), 
  TO_UNSIGNED(419, 12), TO_UNSIGNED(466, 12), 
  TO_UNSIGNED(670, 12), TO_UNSIGNED(712, 12), 
  TO_UNSIGNED(1258, 12), TO_UNSIGNED(1522, 12), 
  TO_UNSIGNED(421, 12), TO_UNSIGNED(468, 12), 
  TO_UNSIGNED(673, 12), TO_UNSIGNED(718, 12), 
  TO_UNSIGNED(1255, 12), TO_UNSIGNED(1546, 12), 
  TO_UNSIGNED(423, 12), TO_UNSIGNED(470, 12), 
  TO_UNSIGNED(676, 12), TO_UNSIGNED(724, 12), 
  TO_UNSIGNED(1264, 12), TO_UNSIGNED(1552, 12), 
  TO_UNSIGNED(425, 12), TO_UNSIGNED(472, 12), 
  TO_UNSIGNED(679, 12), TO_UNSIGNED(730, 12), 
  TO_UNSIGNED(1261, 12), TO_UNSIGNED(1534, 12), 
  TO_UNSIGNED(474, 12), TO_UNSIGNED(522, 12), 
  TO_UNSIGNED(1062, 12), TO_UNSIGNED(1332, 12), 
  TO_UNSIGNED(1631, 12), TO_UNSIGNED(1729, 12), 
  TO_UNSIGNED(476, 12), TO_UNSIGNED(524, 12), 
  TO_UNSIGNED(1068, 12), TO_UNSIGNED(1326, 12), 
  TO_UNSIGNED(1634, 12), TO_UNSIGNED(1723, 12), 
  TO_UNSIGNED(478, 12), TO_UNSIGNED(526, 12), 
  TO_UNSIGNED(1074, 12), TO_UNSIGNED(1350, 12), 
  TO_UNSIGNED(1643, 12), TO_UNSIGNED(1735, 12), 
  TO_UNSIGNED(480, 12), TO_UNSIGNED(528, 12), 
  TO_UNSIGNED(1080, 12), TO_UNSIGNED(1356, 12), 
  TO_UNSIGNED(1640, 12), TO_UNSIGNED(1771, 12), 
  TO_UNSIGNED(482, 12), TO_UNSIGNED(530, 12), 
  TO_UNSIGNED(1086, 12), TO_UNSIGNED(1338, 12), 
  TO_UNSIGNED(1646, 12), TO_UNSIGNED(1777, 12), 
  TO_UNSIGNED(484, 12), TO_UNSIGNED(532, 12), 
  TO_UNSIGNED(1092, 12), TO_UNSIGNED(1344, 12), 
  TO_UNSIGNED(1652, 12), TO_UNSIGNED(1741, 12), 
  TO_UNSIGNED(486, 12), TO_UNSIGNED(534, 12), 
  TO_UNSIGNED(1098, 12), TO_UNSIGNED(1368, 12), 
  TO_UNSIGNED(1649, 12), TO_UNSIGNED(1747, 12), 
  TO_UNSIGNED(488, 12), TO_UNSIGNED(536, 12), 
  TO_UNSIGNED(1104, 12), TO_UNSIGNED(1374, 12), 
  TO_UNSIGNED(1655, 12), TO_UNSIGNED(1753, 12), 
  TO_UNSIGNED(490, 12), TO_UNSIGNED(538, 12), 
  TO_UNSIGNED(1110, 12), TO_UNSIGNED(1362, 12), 
  TO_UNSIGNED(1658, 12), TO_UNSIGNED(1759, 12), 
  TO_UNSIGNED(492, 12), TO_UNSIGNED(540, 12), 
  TO_UNSIGNED(1116, 12), TO_UNSIGNED(1392, 12), 
  TO_UNSIGNED(1661, 12), TO_UNSIGNED(1765, 12), 
  TO_UNSIGNED(494, 12), TO_UNSIGNED(542, 12), 
  TO_UNSIGNED(978, 12), TO_UNSIGNED(1380, 12), 
  TO_UNSIGNED(1664, 12), TO_UNSIGNED(1801, 12), 
  TO_UNSIGNED(496, 12), TO_UNSIGNED(544, 12), 
  TO_UNSIGNED(984, 12), TO_UNSIGNED(1386, 12), 
  TO_UNSIGNED(1667, 12), TO_UNSIGNED(1789, 12), 
  TO_UNSIGNED(130, 12), TO_UNSIGNED(498, 12), 
  TO_UNSIGNED(546, 12), TO_UNSIGNED(990, 12), 
  TO_UNSIGNED(1673, 12), TO_UNSIGNED(1795, 12), 
  TO_UNSIGNED(78, 12), TO_UNSIGNED(500, 12), 
  TO_UNSIGNED(548, 12), TO_UNSIGNED(996, 12), 
  TO_UNSIGNED(1670, 12), TO_UNSIGNED(1807, 12), 
  TO_UNSIGNED(502, 12), TO_UNSIGNED(550, 12), 
  TO_UNSIGNED(1002, 12), TO_UNSIGNED(1272, 12), 
  TO_UNSIGNED(1676, 12), TO_UNSIGNED(1783, 12), 
  TO_UNSIGNED(6, 12), TO_UNSIGNED(504, 12), 
  TO_UNSIGNED(552, 12), TO_UNSIGNED(1008, 12), 
  TO_UNSIGNED(1278, 12), TO_UNSIGNED(1679, 12), 
  TO_UNSIGNED(506, 12), TO_UNSIGNED(554, 12), 
  TO_UNSIGNED(1014, 12), TO_UNSIGNED(1284, 12), 
  TO_UNSIGNED(1682, 12), TO_UNSIGNED(1813, 12), 
  TO_UNSIGNED(136, 12), TO_UNSIGNED(508, 12), 
  TO_UNSIGNED(556, 12), TO_UNSIGNED(1020, 12), 
  TO_UNSIGNED(1266, 12), TO_UNSIGNED(1484, 12), 
  TO_UNSIGNED(510, 12), TO_UNSIGNED(558, 12), 
  TO_UNSIGNED(1026, 12), TO_UNSIGNED(1296, 12), 
  TO_UNSIGNED(1610, 12), TO_UNSIGNED(1687, 12), 
  TO_UNSIGNED(512, 12), TO_UNSIGNED(560, 12), 
  TO_UNSIGNED(1032, 12), TO_UNSIGNED(1290, 12), 
  TO_UNSIGNED(1613, 12), TO_UNSIGNED(1711, 12), 
  TO_UNSIGNED(514, 12), TO_UNSIGNED(562, 12), 
  TO_UNSIGNED(1038, 12), TO_UNSIGNED(1308, 12), 
  TO_UNSIGNED(1622, 12), TO_UNSIGNED(1699, 12), 
  TO_UNSIGNED(516, 12), TO_UNSIGNED(564, 12), 
  TO_UNSIGNED(1044, 12), TO_UNSIGNED(1302, 12), 
  TO_UNSIGNED(1625, 12), TO_UNSIGNED(1705, 12), 
  TO_UNSIGNED(518, 12), TO_UNSIGNED(566, 12), 
  TO_UNSIGNED(1050, 12), TO_UNSIGNED(1314, 12), 
  TO_UNSIGNED(1628, 12), TO_UNSIGNED(1693, 12), 
  TO_UNSIGNED(520, 12), TO_UNSIGNED(568, 12), 
  TO_UNSIGNED(1056, 12), TO_UNSIGNED(1320, 12), 
  TO_UNSIGNED(1637, 12), TO_UNSIGNED(1717, 12), 
  TO_UNSIGNED(523, 12), TO_UNSIGNED(570, 12), 
  TO_UNSIGNED(695, 12), TO_UNSIGNED(877, 12), 
  TO_UNSIGNED(1445, 12), TO_UNSIGNED(1535, 12), 
  TO_UNSIGNED(525, 12), TO_UNSIGNED(572, 12), 
  TO_UNSIGNED(701, 12), TO_UNSIGNED(880, 12), 
  TO_UNSIGNED(1448, 12), TO_UNSIGNED(1541, 12), 
  TO_UNSIGNED(527, 12), TO_UNSIGNED(574, 12), 
  TO_UNSIGNED(707, 12), TO_UNSIGNED(883, 12), 
  TO_UNSIGNED(1451, 12), TO_UNSIGNED(1559, 12), 
  TO_UNSIGNED(529, 12), TO_UNSIGNED(576, 12), 
  TO_UNSIGNED(713, 12), TO_UNSIGNED(886, 12), 
  TO_UNSIGNED(1454, 12), TO_UNSIGNED(1565, 12), 
  TO_UNSIGNED(531, 12), TO_UNSIGNED(578, 12), 
  TO_UNSIGNED(719, 12), TO_UNSIGNED(889, 12), 
  TO_UNSIGNED(1457, 12), TO_UNSIGNED(1577, 12), 
  TO_UNSIGNED(533, 12), TO_UNSIGNED(580, 12), 
  TO_UNSIGNED(725, 12), TO_UNSIGNED(892, 12), 
  TO_UNSIGNED(1463, 12), TO_UNSIGNED(1571, 12), 
  TO_UNSIGNED(535, 12), TO_UNSIGNED(582, 12), 
  TO_UNSIGNED(731, 12), TO_UNSIGNED(895, 12), 
  TO_UNSIGNED(1460, 12), TO_UNSIGNED(1589, 12), 
  TO_UNSIGNED(537, 12), TO_UNSIGNED(584, 12), 
  TO_UNSIGNED(737, 12), TO_UNSIGNED(898, 12), 
  TO_UNSIGNED(1487, 12), TO_UNSIGNED(1583, 12), 
  TO_UNSIGNED(539, 12), TO_UNSIGNED(586, 12), 
  TO_UNSIGNED(743, 12), TO_UNSIGNED(901, 12), 
  TO_UNSIGNED(1601, 12), TO_UNSIGNED(1619, 12), 
  TO_UNSIGNED(541, 12), TO_UNSIGNED(588, 12), 
  TO_UNSIGNED(749, 12), TO_UNSIGNED(904, 12), 
  TO_UNSIGNED(1400, 12), TO_UNSIGNED(1607, 12), 
  TO_UNSIGNED(543, 12), TO_UNSIGNED(590, 12), 
  TO_UNSIGNED(755, 12), TO_UNSIGNED(835, 12), 
  TO_UNSIGNED(1403, 12), TO_UNSIGNED(1595, 12), 
  TO_UNSIGNED(5, 12), TO_UNSIGNED(545, 12), 
  TO_UNSIGNED(592, 12), TO_UNSIGNED(761, 12), 
  TO_UNSIGNED(838, 12), TO_UNSIGNED(1406, 12), 
  TO_UNSIGNED(547, 12), TO_UNSIGNED(594, 12), 
  TO_UNSIGNED(767, 12), TO_UNSIGNED(841, 12), 
  TO_UNSIGNED(1415, 12), TO_UNSIGNED(1481, 12), 
  TO_UNSIGNED(549, 12), TO_UNSIGNED(596, 12), 
  TO_UNSIGNED(773, 12), TO_UNSIGNED(844, 12), 
  TO_UNSIGNED(1418, 12), TO_UNSIGNED(1469, 12), 
  TO_UNSIGNED(551, 12), TO_UNSIGNED(598, 12), 
  TO_UNSIGNED(779, 12), TO_UNSIGNED(847, 12), 
  TO_UNSIGNED(1421, 12), TO_UNSIGNED(1475, 12), 
  TO_UNSIGNED(553, 12), TO_UNSIGNED(600, 12), 
  TO_UNSIGNED(785, 12), TO_UNSIGNED(850, 12), 
  TO_UNSIGNED(1409, 12), TO_UNSIGNED(1499, 12), 
  TO_UNSIGNED(555, 12), TO_UNSIGNED(602, 12), 
  TO_UNSIGNED(791, 12), TO_UNSIGNED(853, 12), 
  TO_UNSIGNED(1412, 12), TO_UNSIGNED(1505, 12), 
  TO_UNSIGNED(557, 12), TO_UNSIGNED(604, 12), 
  TO_UNSIGNED(797, 12), TO_UNSIGNED(856, 12), 
  TO_UNSIGNED(1436, 12), TO_UNSIGNED(1511, 12), 
  TO_UNSIGNED(559, 12), TO_UNSIGNED(606, 12), 
  TO_UNSIGNED(803, 12), TO_UNSIGNED(859, 12), 
  TO_UNSIGNED(1433, 12), TO_UNSIGNED(1493, 12), 
  TO_UNSIGNED(561, 12), TO_UNSIGNED(608, 12), 
  TO_UNSIGNED(809, 12), TO_UNSIGNED(862, 12), 
  TO_UNSIGNED(1424, 12), TO_UNSIGNED(1517, 12), 
  TO_UNSIGNED(563, 12), TO_UNSIGNED(610, 12), 
  TO_UNSIGNED(815, 12), TO_UNSIGNED(865, 12), 
  TO_UNSIGNED(1427, 12), TO_UNSIGNED(1529, 12), 
  TO_UNSIGNED(565, 12), TO_UNSIGNED(612, 12), 
  TO_UNSIGNED(821, 12), TO_UNSIGNED(868, 12), 
  TO_UNSIGNED(1430, 12), TO_UNSIGNED(1523, 12), 
  TO_UNSIGNED(567, 12), TO_UNSIGNED(614, 12), 
  TO_UNSIGNED(827, 12), TO_UNSIGNED(871, 12), 
  TO_UNSIGNED(1439, 12), TO_UNSIGNED(1547, 12), 
  TO_UNSIGNED(569, 12), TO_UNSIGNED(616, 12), 
  TO_UNSIGNED(833, 12), TO_UNSIGNED(874, 12), 
  TO_UNSIGNED(1442, 12), TO_UNSIGNED(1553, 12), 
  TO_UNSIGNED(76, 12), TO_UNSIGNED(571, 12), 
  TO_UNSIGNED(922, 12), TO_UNSIGNED(1105, 12), 
  TO_UNSIGNED(1339, 12), TO_UNSIGNED(1796, 12), 
  TO_UNSIGNED(573, 12), TO_UNSIGNED(925, 12), 
  TO_UNSIGNED(1111, 12), TO_UNSIGNED(1345, 12), 
  TO_UNSIGNED(1615, 12), TO_UNSIGNED(1808, 12), 
  TO_UNSIGNED(575, 12), TO_UNSIGNED(928, 12), 
  TO_UNSIGNED(1117, 12), TO_UNSIGNED(1369, 12), 
  TO_UNSIGNED(1784, 12), TO_UNSIGNED(1820, 12), 
  TO_UNSIGNED(7, 12), TO_UNSIGNED(13, 12), 
  TO_UNSIGNED(577, 12), TO_UNSIGNED(931, 12), 
  TO_UNSIGNED(979, 12), TO_UNSIGNED(1375, 12), 
  TO_UNSIGNED(16, 12), TO_UNSIGNED(579, 12), 
  TO_UNSIGNED(934, 12), TO_UNSIGNED(985, 12), 
  TO_UNSIGNED(1363, 12), TO_UNSIGNED(1814, 12), 
  TO_UNSIGNED(19, 12), TO_UNSIGNED(137, 12), 
  TO_UNSIGNED(581, 12), TO_UNSIGNED(937, 12), 
  TO_UNSIGNED(991, 12), TO_UNSIGNED(1393, 12), 
  TO_UNSIGNED(22, 12), TO_UNSIGNED(583, 12), 
  TO_UNSIGNED(940, 12), TO_UNSIGNED(997, 12), 
  TO_UNSIGNED(1381, 12), TO_UNSIGNED(1688, 12), 
  TO_UNSIGNED(25, 12), TO_UNSIGNED(585, 12), 
  TO_UNSIGNED(943, 12), TO_UNSIGNED(1003, 12), 
  TO_UNSIGNED(1387, 12), TO_UNSIGNED(1712, 12), 
  TO_UNSIGNED(28, 12), TO_UNSIGNED(131, 12), 
  TO_UNSIGNED(587, 12), TO_UNSIGNED(946, 12), 
  TO_UNSIGNED(1009, 12), TO_UNSIGNED(1700, 12), 
  TO_UNSIGNED(31, 12), TO_UNSIGNED(79, 12), 
  TO_UNSIGNED(589, 12), TO_UNSIGNED(949, 12), 
  TO_UNSIGNED(1015, 12), TO_UNSIGNED(1706, 12), 
  TO_UNSIGNED(34, 12), TO_UNSIGNED(591, 12), 
  TO_UNSIGNED(952, 12), TO_UNSIGNED(1021, 12), 
  TO_UNSIGNED(1273, 12), TO_UNSIGNED(1694, 12), 
  TO_UNSIGNED(37, 12), TO_UNSIGNED(593, 12), 
  TO_UNSIGNED(955, 12), TO_UNSIGNED(1027, 12), 
  TO_UNSIGNED(1279, 12), TO_UNSIGNED(1718, 12), 
  TO_UNSIGNED(40, 12), TO_UNSIGNED(595, 12), 
  TO_UNSIGNED(958, 12), TO_UNSIGNED(1033, 12), 
  TO_UNSIGNED(1285, 12), TO_UNSIGNED(1730, 12), 
  TO_UNSIGNED(43, 12), TO_UNSIGNED(597, 12), 
  TO_UNSIGNED(961, 12), TO_UNSIGNED(1039, 12), 
  TO_UNSIGNED(1267, 12), TO_UNSIGNED(1724, 12), 
  TO_UNSIGNED(46, 12), TO_UNSIGNED(599, 12), 
  TO_UNSIGNED(964, 12), TO_UNSIGNED(1045, 12), 
  TO_UNSIGNED(1297, 12), TO_UNSIGNED(1736, 12), 
  TO_UNSIGNED(49, 12), TO_UNSIGNED(601, 12), 
  TO_UNSIGNED(967, 12), TO_UNSIGNED(1051, 12), 
  TO_UNSIGNED(1291, 12), TO_UNSIGNED(1772, 12), 
  TO_UNSIGNED(52, 12), TO_UNSIGNED(603, 12), 
  TO_UNSIGNED(970, 12), TO_UNSIGNED(1057, 12), 
  TO_UNSIGNED(1309, 12), TO_UNSIGNED(1778, 12), 
  TO_UNSIGNED(55, 12), TO_UNSIGNED(605, 12), 
  TO_UNSIGNED(973, 12), TO_UNSIGNED(1063, 12), 
  TO_UNSIGNED(1303, 12), TO_UNSIGNED(1742, 12), 
  TO_UNSIGNED(58, 12), TO_UNSIGNED(607, 12), 
  TO_UNSIGNED(976, 12), TO_UNSIGNED(1069, 12), 
  TO_UNSIGNED(1315, 12), TO_UNSIGNED(1748, 12), 
  TO_UNSIGNED(61, 12), TO_UNSIGNED(609, 12), 
  TO_UNSIGNED(907, 12), TO_UNSIGNED(1075, 12), 
  TO_UNSIGNED(1321, 12), TO_UNSIGNED(1754, 12), 
  TO_UNSIGNED(64, 12), TO_UNSIGNED(611, 12), 
  TO_UNSIGNED(910, 12), TO_UNSIGNED(1081, 12), 
  TO_UNSIGNED(1333, 12), TO_UNSIGNED(1760, 12), 
  TO_UNSIGNED(67, 12), TO_UNSIGNED(613, 12), 
  TO_UNSIGNED(913, 12), TO_UNSIGNED(1087, 12), 
  TO_UNSIGNED(1327, 12), TO_UNSIGNED(1766, 12), 
  TO_UNSIGNED(70, 12), TO_UNSIGNED(615, 12), 
  TO_UNSIGNED(916, 12), TO_UNSIGNED(1093, 12), 
  TO_UNSIGNED(1351, 12), TO_UNSIGNED(1802, 12), 
  TO_UNSIGNED(73, 12), TO_UNSIGNED(617, 12), 
  TO_UNSIGNED(919, 12), TO_UNSIGNED(1099, 12), 
  TO_UNSIGNED(1357, 12), TO_UNSIGNED(1790, 12), 
  TO_UNSIGNED(8, 12), TO_UNSIGNED(132, 12), 
  TO_UNSIGNED(671, 12), TO_UNSIGNED(1028, 12), 
  TO_UNSIGNED(1196, 12), TO_UNSIGNED(1684, 12), 
  TO_UNSIGNED(1685, 12), TO_UNSIGNED(80, 12), 
  TO_UNSIGNED(85, 12), TO_UNSIGNED(674, 12), 
  TO_UNSIGNED(1034, 12), TO_UNSIGNED(1217, 12), 
  TO_UNSIGNED(1815, 12), TO_UNSIGNED(1822, 12), 
  TO_UNSIGNED(87, 12), TO_UNSIGNED(138, 12), 
  TO_UNSIGNED(142, 12), TO_UNSIGNED(677, 12), 
  TO_UNSIGNED(1040, 12), TO_UNSIGNED(1214, 12), 
  TO_UNSIGNED(1274, 12), TO_UNSIGNED(89, 12), 
  TO_UNSIGNED(144, 12), TO_UNSIGNED(680, 12), 
  TO_UNSIGNED(1046, 12), TO_UNSIGNED(1223, 12), 
  TO_UNSIGNED(1280, 12), TO_UNSIGNED(1689, 12), 
  TO_UNSIGNED(91, 12), TO_UNSIGNED(146, 12), 
  TO_UNSIGNED(683, 12), TO_UNSIGNED(1052, 12), 
  TO_UNSIGNED(1226, 12), TO_UNSIGNED(1286, 12), 
  TO_UNSIGNED(1713, 12), TO_UNSIGNED(93, 12), 
  TO_UNSIGNED(148, 12), TO_UNSIGNED(686, 12), 
  TO_UNSIGNED(1058, 12), TO_UNSIGNED(1229, 12), 
  TO_UNSIGNED(1268, 12), TO_UNSIGNED(1701, 12), 
  TO_UNSIGNED(95, 12), TO_UNSIGNED(150, 12), 
  TO_UNSIGNED(689, 12), TO_UNSIGNED(1064, 12), 
  TO_UNSIGNED(1220, 12), TO_UNSIGNED(1298, 12), 
  TO_UNSIGNED(1707, 12), TO_UNSIGNED(97, 12), 
  TO_UNSIGNED(152, 12), TO_UNSIGNED(620, 12), 
  TO_UNSIGNED(1070, 12), TO_UNSIGNED(1235, 12), 
  TO_UNSIGNED(1292, 12), TO_UNSIGNED(1695, 12), 
  TO_UNSIGNED(99, 12), TO_UNSIGNED(154, 12), 
  TO_UNSIGNED(623, 12), TO_UNSIGNED(1076, 12), 
  TO_UNSIGNED(1238, 12), TO_UNSIGNED(1310, 12), 
  TO_UNSIGNED(1719, 12), TO_UNSIGNED(101, 12), 
  TO_UNSIGNED(156, 12), TO_UNSIGNED(626, 12), 
  TO_UNSIGNED(1082, 12), TO_UNSIGNED(1241, 12), 
  TO_UNSIGNED(1304, 12), TO_UNSIGNED(1731, 12), 
  TO_UNSIGNED(103, 12), TO_UNSIGNED(158, 12), 
  TO_UNSIGNED(629, 12), TO_UNSIGNED(1088, 12), 
  TO_UNSIGNED(1232, 12), TO_UNSIGNED(1316, 12), 
  TO_UNSIGNED(1725, 12), TO_UNSIGNED(105, 12), 
  TO_UNSIGNED(160, 12), TO_UNSIGNED(632, 12), 
  TO_UNSIGNED(1094, 12), TO_UNSIGNED(1253, 12), 
  TO_UNSIGNED(1322, 12), TO_UNSIGNED(1737, 12), 
  TO_UNSIGNED(107, 12), TO_UNSIGNED(162, 12), 
  TO_UNSIGNED(635, 12), TO_UNSIGNED(1100, 12), 
  TO_UNSIGNED(1244, 12), TO_UNSIGNED(1334, 12), 
  TO_UNSIGNED(1773, 12), TO_UNSIGNED(109, 12), 
  TO_UNSIGNED(164, 12), TO_UNSIGNED(638, 12), 
  TO_UNSIGNED(1106, 12), TO_UNSIGNED(1247, 12), 
  TO_UNSIGNED(1328, 12), TO_UNSIGNED(1779, 12), 
  TO_UNSIGNED(111, 12), TO_UNSIGNED(166, 12), 
  TO_UNSIGNED(641, 12), TO_UNSIGNED(1112, 12), 
  TO_UNSIGNED(1250, 12), TO_UNSIGNED(1352, 12), 
  TO_UNSIGNED(1743, 12), TO_UNSIGNED(113, 12), 
  TO_UNSIGNED(168, 12), TO_UNSIGNED(644, 12), 
  TO_UNSIGNED(1118, 12), TO_UNSIGNED(1259, 12), 
  TO_UNSIGNED(1358, 12), TO_UNSIGNED(1749, 12), 
  TO_UNSIGNED(115, 12), TO_UNSIGNED(170, 12), 
  TO_UNSIGNED(647, 12), TO_UNSIGNED(980, 12), 
  TO_UNSIGNED(1256, 12), TO_UNSIGNED(1340, 12), 
  TO_UNSIGNED(1755, 12), TO_UNSIGNED(117, 12), 
  TO_UNSIGNED(172, 12), TO_UNSIGNED(650, 12), 
  TO_UNSIGNED(986, 12), TO_UNSIGNED(1265, 12), 
  TO_UNSIGNED(1346, 12), TO_UNSIGNED(1761, 12), 
  TO_UNSIGNED(119, 12), TO_UNSIGNED(174, 12), 
  TO_UNSIGNED(653, 12), TO_UNSIGNED(992, 12), 
  TO_UNSIGNED(1262, 12), TO_UNSIGNED(1370, 12), 
  TO_UNSIGNED(1767, 12), TO_UNSIGNED(121, 12), 
  TO_UNSIGNED(176, 12), TO_UNSIGNED(656, 12), 
  TO_UNSIGNED(998, 12), TO_UNSIGNED(1199, 12), 
  TO_UNSIGNED(1376, 12), TO_UNSIGNED(1803, 12), 
  TO_UNSIGNED(123, 12), TO_UNSIGNED(178, 12), 
  TO_UNSIGNED(659, 12), TO_UNSIGNED(1004, 12), 
  TO_UNSIGNED(1202, 12), TO_UNSIGNED(1364, 12), 
  TO_UNSIGNED(1791, 12), TO_UNSIGNED(125, 12), 
  TO_UNSIGNED(180, 12), TO_UNSIGNED(662, 12), 
  TO_UNSIGNED(1010, 12), TO_UNSIGNED(1205, 12), 
  TO_UNSIGNED(1394, 12), TO_UNSIGNED(1797, 12), 
  TO_UNSIGNED(127, 12), TO_UNSIGNED(182, 12), 
  TO_UNSIGNED(665, 12), TO_UNSIGNED(1016, 12), 
  TO_UNSIGNED(1208, 12), TO_UNSIGNED(1382, 12), 
  TO_UNSIGNED(1809, 12), TO_UNSIGNED(129, 12), 
  TO_UNSIGNED(184, 12), TO_UNSIGNED(668, 12), 
  TO_UNSIGNED(1022, 12), TO_UNSIGNED(1211, 12), 
  TO_UNSIGNED(1388, 12), TO_UNSIGNED(1785, 12), 
  TO_UNSIGNED(187, 12), TO_UNSIGNED(836, 12), 
  TO_UNSIGNED(1083, 12), TO_UNSIGNED(1140, 12), 
  TO_UNSIGNED(1371, 12), TO_UNSIGNED(1686, 12), 
  TO_UNSIGNED(1690, 12), TO_UNSIGNED(189, 12), 
  TO_UNSIGNED(839, 12), TO_UNSIGNED(1089, 12), 
  TO_UNSIGNED(1143, 12), TO_UNSIGNED(1377, 12), 
  TO_UNSIGNED(1714, 12), TO_UNSIGNED(1823, 12), 
  TO_UNSIGNED(143, 12), TO_UNSIGNED(191, 12), 
  TO_UNSIGNED(842, 12), TO_UNSIGNED(1095, 12), 
  TO_UNSIGNED(1146, 12), TO_UNSIGNED(1365, 12), 
  TO_UNSIGNED(1702, 12), TO_UNSIGNED(145, 12), 
  TO_UNSIGNED(193, 12), TO_UNSIGNED(845, 12), 
  TO_UNSIGNED(1101, 12), TO_UNSIGNED(1149, 12), 
  TO_UNSIGNED(1395, 12), TO_UNSIGNED(1708, 12), 
  TO_UNSIGNED(147, 12), TO_UNSIGNED(195, 12), 
  TO_UNSIGNED(848, 12), TO_UNSIGNED(1107, 12), 
  TO_UNSIGNED(1152, 12), TO_UNSIGNED(1383, 12), 
  TO_UNSIGNED(1696, 12), TO_UNSIGNED(149, 12), 
  TO_UNSIGNED(197, 12), TO_UNSIGNED(851, 12), 
  TO_UNSIGNED(1113, 12), TO_UNSIGNED(1155, 12), 
  TO_UNSIGNED(1389, 12), TO_UNSIGNED(1720, 12), 
  TO_UNSIGNED(133, 12), TO_UNSIGNED(151, 12), 
  TO_UNSIGNED(199, 12), TO_UNSIGNED(854, 12), 
  TO_UNSIGNED(1119, 12), TO_UNSIGNED(1158, 12), 
  TO_UNSIGNED(1732, 12), TO_UNSIGNED(81, 12), 
  TO_UNSIGNED(153, 12), TO_UNSIGNED(201, 12), 
  TO_UNSIGNED(857, 12), TO_UNSIGNED(981, 12), 
  TO_UNSIGNED(1161, 12), TO_UNSIGNED(1726, 12), 
  TO_UNSIGNED(155, 12), TO_UNSIGNED(203, 12), 
  TO_UNSIGNED(860, 12), TO_UNSIGNED(987, 12), 
  TO_UNSIGNED(1164, 12), TO_UNSIGNED(1275, 12), 
  TO_UNSIGNED(1738, 12), TO_UNSIGNED(157, 12), 
  TO_UNSIGNED(205, 12), TO_UNSIGNED(863, 12), 
  TO_UNSIGNED(993, 12), TO_UNSIGNED(1167, 12), 
  TO_UNSIGNED(1281, 12), TO_UNSIGNED(1774, 12), 
  TO_UNSIGNED(159, 12), TO_UNSIGNED(207, 12), 
  TO_UNSIGNED(866, 12), TO_UNSIGNED(999, 12), 
  TO_UNSIGNED(1170, 12), TO_UNSIGNED(1287, 12), 
  TO_UNSIGNED(1780, 12), TO_UNSIGNED(161, 12), 
  TO_UNSIGNED(209, 12), TO_UNSIGNED(869, 12), 
  TO_UNSIGNED(1005, 12), TO_UNSIGNED(1173, 12), 
  TO_UNSIGNED(1269, 12), TO_UNSIGNED(1744, 12), 
  TO_UNSIGNED(163, 12), TO_UNSIGNED(211, 12), 
  TO_UNSIGNED(872, 12), TO_UNSIGNED(1011, 12), 
  TO_UNSIGNED(1176, 12), TO_UNSIGNED(1299, 12), 
  TO_UNSIGNED(1750, 12), TO_UNSIGNED(165, 12), 
  TO_UNSIGNED(213, 12), TO_UNSIGNED(875, 12), 
  TO_UNSIGNED(1017, 12), TO_UNSIGNED(1179, 12), 
  TO_UNSIGNED(1293, 12), TO_UNSIGNED(1756, 12), 
  TO_UNSIGNED(167, 12), TO_UNSIGNED(215, 12), 
  TO_UNSIGNED(878, 12), TO_UNSIGNED(1023, 12), 
  TO_UNSIGNED(1182, 12), TO_UNSIGNED(1311, 12), 
  TO_UNSIGNED(1762, 12), TO_UNSIGNED(169, 12), 
  TO_UNSIGNED(217, 12), TO_UNSIGNED(881, 12), 
  TO_UNSIGNED(1029, 12), TO_UNSIGNED(1185, 12), 
  TO_UNSIGNED(1305, 12), TO_UNSIGNED(1768, 12), 
  TO_UNSIGNED(171, 12), TO_UNSIGNED(219, 12), 
  TO_UNSIGNED(884, 12), TO_UNSIGNED(1035, 12), 
  TO_UNSIGNED(1188, 12), TO_UNSIGNED(1317, 12), 
  TO_UNSIGNED(1804, 12), TO_UNSIGNED(173, 12), 
  TO_UNSIGNED(221, 12), TO_UNSIGNED(887, 12), 
  TO_UNSIGNED(1041, 12), TO_UNSIGNED(1191, 12), 
  TO_UNSIGNED(1323, 12), TO_UNSIGNED(1792, 12), 
  TO_UNSIGNED(175, 12), TO_UNSIGNED(223, 12), 
  TO_UNSIGNED(890, 12), TO_UNSIGNED(1047, 12), 
  TO_UNSIGNED(1122, 12), TO_UNSIGNED(1335, 12), 
  TO_UNSIGNED(1798, 12), TO_UNSIGNED(177, 12), 
  TO_UNSIGNED(225, 12), TO_UNSIGNED(893, 12), 
  TO_UNSIGNED(1053, 12), TO_UNSIGNED(1125, 12), 
  TO_UNSIGNED(1329, 12), TO_UNSIGNED(1810, 12), 
  TO_UNSIGNED(179, 12), TO_UNSIGNED(227, 12), 
  TO_UNSIGNED(896, 12), TO_UNSIGNED(1059, 12), 
  TO_UNSIGNED(1128, 12), TO_UNSIGNED(1353, 12), 
  TO_UNSIGNED(1786, 12), TO_UNSIGNED(9, 12), 
  TO_UNSIGNED(181, 12), TO_UNSIGNED(229, 12), 
  TO_UNSIGNED(899, 12), TO_UNSIGNED(1065, 12), 
  TO_UNSIGNED(1131, 12), TO_UNSIGNED(1359, 12), 
  TO_UNSIGNED(183, 12), TO_UNSIGNED(231, 12), 
  TO_UNSIGNED(902, 12), TO_UNSIGNED(1071, 12), 
  TO_UNSIGNED(1134, 12), TO_UNSIGNED(1341, 12), 
  TO_UNSIGNED(1816, 12), TO_UNSIGNED(139, 12), 
  TO_UNSIGNED(185, 12), TO_UNSIGNED(233, 12), 
  TO_UNSIGNED(905, 12), TO_UNSIGNED(1077, 12), 
  TO_UNSIGNED(1137, 12), TO_UNSIGNED(1347, 12), 
  TO_UNSIGNED(283, 12), TO_UNSIGNED(331, 12), 
  TO_UNSIGNED(1000, 12), TO_UNSIGNED(1123, 12), 
  TO_UNSIGNED(1300, 12), TO_UNSIGNED(1616, 12), 
  TO_UNSIGNED(1721, 12), TO_UNSIGNED(285, 12), 
  TO_UNSIGNED(333, 12), TO_UNSIGNED(1006, 12), 
  TO_UNSIGNED(1126, 12), TO_UNSIGNED(1294, 12), 
  TO_UNSIGNED(1733, 12), TO_UNSIGNED(1821, 12), 
  TO_UNSIGNED(14, 12), TO_UNSIGNED(287, 12), 
  TO_UNSIGNED(335, 12), TO_UNSIGNED(1012, 12), 
  TO_UNSIGNED(1129, 12), TO_UNSIGNED(1312, 12), 
  TO_UNSIGNED(1727, 12), TO_UNSIGNED(17, 12), 
  TO_UNSIGNED(289, 12), TO_UNSIGNED(337, 12), 
  TO_UNSIGNED(1018, 12), TO_UNSIGNED(1132, 12), 
  TO_UNSIGNED(1306, 12), TO_UNSIGNED(1739, 12), 
  TO_UNSIGNED(20, 12), TO_UNSIGNED(291, 12), 
  TO_UNSIGNED(339, 12), TO_UNSIGNED(1024, 12), 
  TO_UNSIGNED(1135, 12), TO_UNSIGNED(1318, 12), 
  TO_UNSIGNED(1775, 12), TO_UNSIGNED(23, 12), 
  TO_UNSIGNED(293, 12), TO_UNSIGNED(341, 12), 
  TO_UNSIGNED(1030, 12), TO_UNSIGNED(1138, 12), 
  TO_UNSIGNED(1324, 12), TO_UNSIGNED(1781, 12), 
  TO_UNSIGNED(26, 12), TO_UNSIGNED(295, 12), 
  TO_UNSIGNED(343, 12), TO_UNSIGNED(1036, 12), 
  TO_UNSIGNED(1141, 12), TO_UNSIGNED(1336, 12), 
  TO_UNSIGNED(1745, 12), TO_UNSIGNED(29, 12), 
  TO_UNSIGNED(297, 12), TO_UNSIGNED(345, 12), 
  TO_UNSIGNED(1042, 12), TO_UNSIGNED(1144, 12), 
  TO_UNSIGNED(1330, 12), TO_UNSIGNED(1751, 12), 
  TO_UNSIGNED(32, 12), TO_UNSIGNED(299, 12), 
  TO_UNSIGNED(347, 12), TO_UNSIGNED(1048, 12), 
  TO_UNSIGNED(1147, 12), TO_UNSIGNED(1354, 12), 
  TO_UNSIGNED(1757, 12), TO_UNSIGNED(35, 12), 
  TO_UNSIGNED(301, 12), TO_UNSIGNED(349, 12), 
  TO_UNSIGNED(1054, 12), TO_UNSIGNED(1150, 12), 
  TO_UNSIGNED(1360, 12), TO_UNSIGNED(1763, 12), 
  TO_UNSIGNED(38, 12), TO_UNSIGNED(303, 12), 
  TO_UNSIGNED(351, 12), TO_UNSIGNED(1060, 12), 
  TO_UNSIGNED(1153, 12), TO_UNSIGNED(1342, 12), 
  TO_UNSIGNED(1769, 12), TO_UNSIGNED(41, 12), 
  TO_UNSIGNED(305, 12), TO_UNSIGNED(353, 12), 
  TO_UNSIGNED(1066, 12), TO_UNSIGNED(1156, 12), 
  TO_UNSIGNED(1348, 12), TO_UNSIGNED(1805, 12), 
  TO_UNSIGNED(44, 12), TO_UNSIGNED(307, 12), 
  TO_UNSIGNED(355, 12), TO_UNSIGNED(1072, 12), 
  TO_UNSIGNED(1159, 12), TO_UNSIGNED(1372, 12), 
  TO_UNSIGNED(1793, 12), TO_UNSIGNED(47, 12), 
  TO_UNSIGNED(309, 12), TO_UNSIGNED(357, 12), 
  TO_UNSIGNED(1078, 12), TO_UNSIGNED(1162, 12), 
  TO_UNSIGNED(1378, 12), TO_UNSIGNED(1799, 12), 
  TO_UNSIGNED(50, 12), TO_UNSIGNED(311, 12), 
  TO_UNSIGNED(359, 12), TO_UNSIGNED(1084, 12), 
  TO_UNSIGNED(1165, 12), TO_UNSIGNED(1366, 12), 
  TO_UNSIGNED(1811, 12), TO_UNSIGNED(53, 12), 
  TO_UNSIGNED(313, 12), TO_UNSIGNED(361, 12), 
  TO_UNSIGNED(1090, 12), TO_UNSIGNED(1168, 12), 
  TO_UNSIGNED(1396, 12), TO_UNSIGNED(1787, 12), 
  TO_UNSIGNED(10, 12), TO_UNSIGNED(56, 12), 
  TO_UNSIGNED(315, 12), TO_UNSIGNED(363, 12), 
  TO_UNSIGNED(1096, 12), TO_UNSIGNED(1171, 12), 
  TO_UNSIGNED(1384, 12), TO_UNSIGNED(59, 12), 
  TO_UNSIGNED(317, 12), TO_UNSIGNED(365, 12), 
  TO_UNSIGNED(1102, 12), TO_UNSIGNED(1174, 12), 
  TO_UNSIGNED(1390, 12), TO_UNSIGNED(1817, 12), 
  TO_UNSIGNED(62, 12), TO_UNSIGNED(134, 12), 
  TO_UNSIGNED(140, 12), TO_UNSIGNED(319, 12), 
  TO_UNSIGNED(367, 12), TO_UNSIGNED(1108, 12), 
  TO_UNSIGNED(1177, 12), TO_UNSIGNED(65, 12), 
  TO_UNSIGNED(82, 12), TO_UNSIGNED(321, 12), 
  TO_UNSIGNED(369, 12), TO_UNSIGNED(1114, 12), 
  TO_UNSIGNED(1180, 12), TO_UNSIGNED(1691, 12), 
  TO_UNSIGNED(68, 12), TO_UNSIGNED(323, 12), 
  TO_UNSIGNED(371, 12), TO_UNSIGNED(1120, 12), 
  TO_UNSIGNED(1183, 12), TO_UNSIGNED(1276, 12), 
  TO_UNSIGNED(1715, 12), TO_UNSIGNED(71, 12), 
  TO_UNSIGNED(325, 12), TO_UNSIGNED(373, 12), 
  TO_UNSIGNED(982, 12), TO_UNSIGNED(1186, 12), 
  TO_UNSIGNED(1282, 12), TO_UNSIGNED(1703, 12), 
  TO_UNSIGNED(74, 12), TO_UNSIGNED(327, 12), 
  TO_UNSIGNED(375, 12), TO_UNSIGNED(988, 12), 
  TO_UNSIGNED(1189, 12), TO_UNSIGNED(1288, 12), 
  TO_UNSIGNED(1709, 12), TO_UNSIGNED(77, 12), 
  TO_UNSIGNED(329, 12), TO_UNSIGNED(377, 12), 
  TO_UNSIGNED(994, 12), TO_UNSIGNED(1192, 12), 
  TO_UNSIGNED(1270, 12), TO_UNSIGNED(1697, 12), 
  TO_UNSIGNED(427, 12), TO_UNSIGNED(475, 12), 
  TO_UNSIGNED(944, 12), TO_UNSIGNED(1025, 12), 
  TO_UNSIGNED(1169, 12), TO_UNSIGNED(1343, 12), 
  TO_UNSIGNED(1752, 12), TO_UNSIGNED(429, 12), 
  TO_UNSIGNED(477, 12), TO_UNSIGNED(947, 12), 
  TO_UNSIGNED(1031, 12), TO_UNSIGNED(1172, 12), 
  TO_UNSIGNED(1349, 12), TO_UNSIGNED(1758, 12), 
  TO_UNSIGNED(431, 12), TO_UNSIGNED(479, 12), 
  TO_UNSIGNED(950, 12), TO_UNSIGNED(1037, 12), 
  TO_UNSIGNED(1175, 12), TO_UNSIGNED(1373, 12), 
  TO_UNSIGNED(1764, 12), TO_UNSIGNED(433, 12), 
  TO_UNSIGNED(481, 12), TO_UNSIGNED(953, 12), 
  TO_UNSIGNED(1043, 12), TO_UNSIGNED(1178, 12), 
  TO_UNSIGNED(1379, 12), TO_UNSIGNED(1770, 12), 
  TO_UNSIGNED(435, 12), TO_UNSIGNED(483, 12), 
  TO_UNSIGNED(956, 12), TO_UNSIGNED(1049, 12), 
  TO_UNSIGNED(1181, 12), TO_UNSIGNED(1367, 12), 
  TO_UNSIGNED(1806, 12), TO_UNSIGNED(437, 12), 
  TO_UNSIGNED(485, 12), TO_UNSIGNED(959, 12), 
  TO_UNSIGNED(1055, 12), TO_UNSIGNED(1184, 12), 
  TO_UNSIGNED(1397, 12), TO_UNSIGNED(1794, 12), 
  TO_UNSIGNED(439, 12), TO_UNSIGNED(487, 12), 
  TO_UNSIGNED(962, 12), TO_UNSIGNED(1061, 12), 
  TO_UNSIGNED(1187, 12), TO_UNSIGNED(1385, 12), 
  TO_UNSIGNED(1800, 12), TO_UNSIGNED(441, 12), 
  TO_UNSIGNED(489, 12), TO_UNSIGNED(965, 12), 
  TO_UNSIGNED(1067, 12), TO_UNSIGNED(1190, 12), 
  TO_UNSIGNED(1391, 12), TO_UNSIGNED(1812, 12), 
  TO_UNSIGNED(135, 12), TO_UNSIGNED(443, 12), 
  TO_UNSIGNED(491, 12), TO_UNSIGNED(968, 12), 
  TO_UNSIGNED(1073, 12), TO_UNSIGNED(1193, 12), 
  TO_UNSIGNED(1788, 12), TO_UNSIGNED(11, 12), 
  TO_UNSIGNED(83, 12), TO_UNSIGNED(445, 12), 
  TO_UNSIGNED(493, 12), TO_UNSIGNED(971, 12), 
  TO_UNSIGNED(1079, 12), TO_UNSIGNED(1124, 12), 
  TO_UNSIGNED(447, 12), TO_UNSIGNED(495, 12), 
  TO_UNSIGNED(974, 12), TO_UNSIGNED(1085, 12), 
  TO_UNSIGNED(1127, 12), TO_UNSIGNED(1277, 12), 
  TO_UNSIGNED(1818, 12), TO_UNSIGNED(141, 12), 
  TO_UNSIGNED(449, 12), TO_UNSIGNED(497, 12), 
  TO_UNSIGNED(977, 12), TO_UNSIGNED(1091, 12), 
  TO_UNSIGNED(1130, 12), TO_UNSIGNED(1283, 12), 
  TO_UNSIGNED(451, 12), TO_UNSIGNED(499, 12), 
  TO_UNSIGNED(908, 12), TO_UNSIGNED(1097, 12), 
  TO_UNSIGNED(1133, 12), TO_UNSIGNED(1289, 12), 
  TO_UNSIGNED(1692, 12), TO_UNSIGNED(453, 12), 
  TO_UNSIGNED(501, 12), TO_UNSIGNED(911, 12), 
  TO_UNSIGNED(1103, 12), TO_UNSIGNED(1136, 12), 
  TO_UNSIGNED(1271, 12), TO_UNSIGNED(1716, 12), 
  TO_UNSIGNED(455, 12), TO_UNSIGNED(503, 12), 
  TO_UNSIGNED(914, 12), TO_UNSIGNED(1109, 12), 
  TO_UNSIGNED(1139, 12), TO_UNSIGNED(1301, 12), 
  TO_UNSIGNED(1704, 12), TO_UNSIGNED(457, 12), 
  TO_UNSIGNED(505, 12), TO_UNSIGNED(917, 12), 
  TO_UNSIGNED(1115, 12), TO_UNSIGNED(1142, 12), 
  TO_UNSIGNED(1295, 12), TO_UNSIGNED(1710, 12), 
  TO_UNSIGNED(459, 12), TO_UNSIGNED(507, 12), 
  TO_UNSIGNED(920, 12), TO_UNSIGNED(1121, 12), 
  TO_UNSIGNED(1145, 12), TO_UNSIGNED(1313, 12), 
  TO_UNSIGNED(1698, 12), TO_UNSIGNED(461, 12), 
  TO_UNSIGNED(509, 12), TO_UNSIGNED(923, 12), 
  TO_UNSIGNED(983, 12), TO_UNSIGNED(1148, 12), 
  TO_UNSIGNED(1307, 12), TO_UNSIGNED(1722, 12), 
  TO_UNSIGNED(463, 12), TO_UNSIGNED(511, 12), 
  TO_UNSIGNED(926, 12), TO_UNSIGNED(989, 12), 
  TO_UNSIGNED(1151, 12), TO_UNSIGNED(1319, 12), 
  TO_UNSIGNED(1734, 12), TO_UNSIGNED(465, 12), 
  TO_UNSIGNED(513, 12), TO_UNSIGNED(929, 12), 
  TO_UNSIGNED(995, 12), TO_UNSIGNED(1154, 12), 
  TO_UNSIGNED(1325, 12), TO_UNSIGNED(1728, 12), 
  TO_UNSIGNED(467, 12), TO_UNSIGNED(515, 12), 
  TO_UNSIGNED(932, 12), TO_UNSIGNED(1001, 12), 
  TO_UNSIGNED(1157, 12), TO_UNSIGNED(1337, 12), 
  TO_UNSIGNED(1740, 12), TO_UNSIGNED(469, 12), 
  TO_UNSIGNED(517, 12), TO_UNSIGNED(935, 12), 
  TO_UNSIGNED(1007, 12), TO_UNSIGNED(1160, 12), 
  TO_UNSIGNED(1331, 12), TO_UNSIGNED(1776, 12), 
  TO_UNSIGNED(471, 12), TO_UNSIGNED(519, 12), 
  TO_UNSIGNED(938, 12), TO_UNSIGNED(1013, 12), 
  TO_UNSIGNED(1163, 12), TO_UNSIGNED(1355, 12), 
  TO_UNSIGNED(1782, 12), TO_UNSIGNED(473, 12), 
  TO_UNSIGNED(521, 12), TO_UNSIGNED(941, 12), 
  TO_UNSIGNED(1019, 12), TO_UNSIGNED(1166, 12), 
  TO_UNSIGNED(1361, 12), TO_UNSIGNED(1746, 12)
);                        

	SIGNAL READ_C  : UNSIGNED(11 downto 0);
	SIGNAL WRITE_C : UNSIGNED(11 downto 0);
	SIGNAL ROM_ADR : UNSIGNED(11 downto 0);

BEGIN

	-------------------------------------------------------------------------
	-- synthesis translate_off 
  	PROCESS
  	BEGIN
    	WAIT FOR 1 ns;
		--printmsg("(IMS) Q16_8_IndexLUT : ALLOCATION OK !");
    	WAIT;
  	END PROCESS;
	-- synthesis translate_on 
	-------------------------------------------------------------------------

	--
	--
	--
	process(clock, reset)
		VARIABLE TEMP : UNSIGNED(11 downto 0);
	begin
		if reset = '0' then
			WRITE_C <= TO_UNSIGNED(0, 12);
		elsif clock'event and clock = '1' then
			if write_en = '1' then
				TEMP := WRITE_C + TO_UNSIGNED(1, 12);
				IF TEMP = 1824 THEN
					TEMP := TO_UNSIGNED(0, 12);
				END IF;
				WRITE_C <= TEMP;
			else
				WRITE_C <= WRITE_C;
			end if;
			WE_BIS <= write_en;
			IN_BIS <= INPUT_1;
		end if;
	end process;


	--
	--
	--
	process(clock, reset)
		VARIABLE TEMP : UNSIGNED(11 downto 0);
	begin
		if reset = '0' then
			READ_C <= TO_UNSIGNED(0, 12);
		elsif clock'event and clock = '1' then
			if read_en = '1' then
				TEMP := READ_C + TO_UNSIGNED(1, 12);
				IF TEMP = 1824 THEN
					TEMP := TO_UNSIGNED(0, 12);
				END IF;
				READ_C <= TEMP;
			else
				READ_C <= READ_C;
			end if;
		end if;
	end process;


	--
	--
	--
	process(clock)
		VARIABLE ADR : INTEGER RANGE 0 to 1823;
		VARIABLE POS : INTEGER RANGE 0 to 1823;
	begin
		if clock'event and clock = '1' then
			ADR     := to_integer( WRITE_C );
			ROM_ADR <= ROM( ADR );
		end if;
	end process;


	--
	--
	--
	process(clock)
	begin
		if clock'event and clock = '1' then
			if WE_BIS = '1' then
				RAM( to_integer( ROM_ADR ) ) <= IN_BIS;
			end if;
			OUTPUT_1 <= RAM( to_integer(READ_C) );
		end if;
	end process;

END cRAM;
