--	ADDER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY ADD_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

architecture behavior of ADD_Dynamic is
  -- MAXIMUM FUNCTION TO COMPUTE THE INTERNAL DATA SIZE
  FUNCTION maximum (left, right : NATURAL) return NATURAL IS
  BEGIN  -- function max
    IF LEFT > RIGHT THEN RETURN LEFT;
    ELSE RETURN RIGHT;
    END IF;
  END FUNCTION maximum;

BEGIN
	PROCESS (INPUT_1, INPUT_2)
		CONSTANT SIZI  : NATURAL := maximum(INPUT_1_WIDTH, INPUT_2_WIDTH);
		CONSTANT SIZE  : NATURAL := maximum(SIZI, OUTPUT_1_WIDTH);
		VARIABLE Stmp  : SIGNED  (SIZE-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED(SIZE-1 DOWNTO 0);
	BEGIN
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED( INPUT_1 ) + UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH);

			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		ELSE
			Stmp     := RESIZE( SIGNED( INPUT_1 ) + SIGNED( INPUT_2 ), OUTPUT_1_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		END IF;
	END PROCESS;
END;


--	SUBSTRACTOR COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY SUB_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :IN  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

ARCHITECTURE behavior OF SUB_Dynamic IS

  -- MAXIMUM FUNCTION TO COMPUTE THE INTERNAL DATA SIZE
  FUNCTION maximum (left, right : NATURAL) return NATURAL IS
  BEGIN  -- function max
    IF LEFT > RIGHT THEN RETURN LEFT;
    ELSE RETURN RIGHT;
    END IF;
  END FUNCTION maximum;

BEGIN
	PROCESS (INPUT_1, INPUT_2)
		CONSTANT SIZI  : NATURAL := maximum(INPUT_1_WIDTH, INPUT_2_WIDTH);
		CONSTANT SIZE  : NATURAL := maximum(SIZI, OUTPUT_1_WIDTH);
		VARIABLE Stmp  : SIGNED  (SIZE-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED(SIZE-1 DOWNTO 0);
	BEGIN
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED( INPUT_1 ) - UNSIGNED( INPUT_2 ), OUTPUT_1_WIDTH);

			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );

		ELSE

			Stmp     := RESIZE( SIGNED( INPUT_1 ) - SIGNED( INPUT_2 ), OUTPUT_1_WIDTH);

			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );

		END IF;
	END PROCESS;
END;




--	MULTIPLIER COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

entity MUL_Dynamic is
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	INPUT_2_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  port ( 
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		INPUT_2  :in  STD_LOGIC_VECTOR(INPUT_2_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
end;

architecture behavior of MUL_Dynamic is
  -- MAXIMUM FUNCTION TO COMPUTE THE INTERNAL DATA SIZE

  FUNCTION maximum (left, right : NATURAL) return NATURAL IS

  BEGIN  -- function max

    IF LEFT > RIGHT THEN RETURN LEFT;

    ELSE RETURN RIGHT;

    END IF;

  END FUNCTION maximum;



BEGIN

	process (INPUT_1, INPUT_2)
		VARIABLE Stmp  : SIGNED  ((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED((INPUT_1_WIDTH+INPUT_2_WIDTH)-1 DOWNTO 0);
	begin
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED( INPUT_1 ) * UNSIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);

			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );

		ELSE

			Stmp     := RESIZE( SIGNED( INPUT_1 ) * SIGNED( INPUT_2 ), INPUT_1_WIDTH+INPUT_2_WIDTH);

			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );

		END IF;
	end process;
end;


--	SQUARE COMPONENT WITH VARIABLE INPUTS AND OUTPUT BITWIDTH
--	DEVELOPPED FOR THE GRAPHLAB TOOL BY BERTRAND LE GAL
--	IMS LABORATORY -  UMR-CNRS 5218
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

entity SQR_Dynamic is
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  port (
		INPUT_1  :in  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :out STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
end;

architecture behavior of SQR_Dynamic is
begin
	process (INPUT_1)
		VARIABLE Stmp  : SIGNED  ((INPUT_1_WIDTH+INPUT_1_WIDTH)-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED((INPUT_1_WIDTH+INPUT_1_WIDTH)-1 DOWNTO 0);
	begin
		IF C_SIGNED = 0 THEN
			UStmp    := UNSIGNED( INPUT_1 ) * UNSIGNED( INPUT_1 );
			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		ELSE
			Stmp     := SIGNED( INPUT_1 ) * SIGNED( INPUT_1 );
			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		END IF;
	end process;
end;



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;

ENTITY ABS_Dynamic IS
  GENERIC(
      	C_SIGNED          : NATURAL := 0;
      	INPUT_1_WIDTH     : NATURAL := 8;
      	OUTPUT_1_WIDTH    : NATURAL := 8
  	  );
  PORT ( 
		INPUT_1  :IN  STD_LOGIC_VECTOR(INPUT_1_WIDTH-1  DOWNTO 0);
		OUTPUT_1 :OUT STD_LOGIC_VECTOR(OUTPUT_1_WIDTH-1 DOWNTO 0)
		);
END;

architecture behavior of ABS_Dynamic is
  -- MAXIMUM FUNCTION TO COMPUTE THE INTERNAL DATA SIZE
  FUNCTION minimum (left, right : NATURAL) return NATURAL IS
  BEGIN  -- function max
    IF LEFT < RIGHT THEN RETURN LEFT;
    ELSE RETURN RIGHT;
    END IF;
  END FUNCTION minimum;

BEGIN
	PROCESS (INPUT_1)
		CONSTANT SIZE  : NATURAL := minimum(INPUT_1_WIDTH, OUTPUT_1_WIDTH);
		VARIABLE Stmp  : SIGNED  (SIZE-1 DOWNTO 0);
		VARIABLE UStmp : UNSIGNED(SIZE-1 DOWNTO 0);
	BEGIN
		IF C_SIGNED = 0 THEN
			UStmp    := RESIZE( UNSIGNED(INPUT_1), OUTPUT_1_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( UStmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		ELSE
			Stmp     := RESIZE( abs(SIGNED( INPUT_1 )), OUTPUT_1_WIDTH);
			OUTPUT_1 <= STD_LOGIC_VECTOR( Stmp(OUTPUT_1_WIDTH-1 DOWNTO 0) );
		END IF;
	END PROCESS;
END;
