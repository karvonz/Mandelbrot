library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library WORK;
use WORK.CONSTANTS.ALL;
use WORK.FUNCTIONS.ALL;

entity Colorgen is
    Port ( iters : in STD_LOGIC_VECTOR (ITER_RANGE-1 downto 0);
			  itermax : in STD_LOGIC_VECTOR (ITER_RANGE-1 downto 0);
           color : out STD_LOGIC_VECTOR (bit_per_pixel-1 downto 0));
end Colorgen;


architecture Behavioral of Colorgen is
	type  rom_type is array (0 to ITER_MAX-1) of std_logic_vector (bit_per_pixel-1 downto 0);
	constant color_scheme : rom_type := (
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000001",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000010",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000011",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000100",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000101",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000110",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000000111",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001000",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001001",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001010",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001011",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001100",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001101",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001110",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000001111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000011111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000101111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000000111111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001001111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001011111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001101111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000001111111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010001111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010011111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010101111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000010111111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011001111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011011111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011101111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111111",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111110",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111101",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111100",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111011",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111010",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111001",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011111000",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110111",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110110",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110101",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110100",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110011",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110010",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110001",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000011110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"000111110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001011110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"001111110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010011110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"010111110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011011110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"011111110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100011110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"100111110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101011110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"101111110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110011110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"110111110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111011110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"111111110000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000"
);

begin
process(iters, itermax)
begin
	if (iters = itermax) then
		color<= (others=>'0');
	else
		color <= color_scheme(to_integer(unsigned(iters)));
	end if;
end process;end Behavioral;


--Cut and paste following lines into Shared.vhd.
--	constant ITER_MAX : integer := 4095;
--	constant ITER_RANGE : integer := 12;
