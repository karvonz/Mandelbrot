library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library WORK;
use WORK.CONSTANTS.ALL;
use WORK.FUNCTIONS.ALL;

entity Colorgen is
    Port ( iter : in STD_LOGIC_VECTOR (11 downto 0);
	 VGA_red      : out std_logic_vector(3 downto 0);   -- red output
       VGA_green    : out std_logic_vector(3 downto 0);   -- green output
       VGA_blue     : out std_logic_vector(3 downto 0));   -- blue output
end Colorgen;


architecture Behavioral of Colorgen is -- TODO : Am�liorer colorgen (comparaison OpenGL)
	
	
	
	type  rom_type is array (0 to 4095) of std_logic_vector (bit_per_pixel-1 downto 0);
	constant color_scheme : rom_type := (
		x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"001", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"002", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"003", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"004", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"005", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"006", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"007", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"017", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"018", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"019", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02A", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"02B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03B", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"03C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04C", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"04D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"05D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"06D", 
x"16D", 
x"16D", 
x"16D", 
x"16D", 
x"16D", 
x"16D", 
x"16D", 
x"16D", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"16E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"17E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"18E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"19E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"29E", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AE", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2AD", 
x"2BD", 
x"2BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3BD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"3CD", 
x"4CD", 
x"4CD", 
x"4CD", 
x"4CD", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4CC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"4DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DC", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5DB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"5EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EB", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"6EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7EA", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"7E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E9", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"8E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E8", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"9E7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE7", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"AE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE6", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"BE5", 
x"CE5", 
x"CE5", 
x"CE5", 
x"CE5", 
x"CE5", 
x"CE5", 
x"CE5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD5", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"CD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DD4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC4", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"DC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EC3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB3", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EB2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"EA2", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"E92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F92", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F91", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F81", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"F71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E71", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E61", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E60", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E50", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"E40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D40", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"D30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C30", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"C20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"B20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A20", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"A10", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"910", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"810", 
x"800", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"700", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"600", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"500", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"400", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"300", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"200", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"100", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000", 
x"000"
);

begin
process(iter)
begin
	--color <= not iters;
	
	           VGA_red   <= color_scheme(to_integer(unsigned(iter)))(11 downto 8);
               VGA_green <= color_scheme(to_integer(unsigned(iter)))( 7 downto 4);
               VGA_blue  <= color_scheme(to_integer(unsigned(iter)))( 3 downto 0);

end process;

end Behavioral;


--Cut and paste following lines into Shared.vhd.
--	constant ITER_MAX : integer := 4095;
--	constant ITER_RANGE : integer := 12;
